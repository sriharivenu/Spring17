
module fifo_DW01_mux_any_256_4_16_1 ( A, SEL, MUX );
input  [255:0] A;
input  [3:0] SEL;
output [15:0] MUX;
    wire \tmp[3][136] , \tmp[3][14] , \tmp[3][132] , \tmp[3][10] , 
        \tmp[3][139] , \tmp[3][130] , \tmp[3][129] , \tmp[3][12] , 
        \tmp[3][134] , \tmp[3][1] , \tmp[3][8] , \tmp[3][141] , \tmp[3][5] , 
        \tmp[3][7] , \tmp[3][143] , \tmp[3][3] , \tmp[3][142] , \tmp[3][2] , 
        \tmp[3][6] , \tmp[3][4] , \tmp[3][0] , \tmp[3][9] , \tmp[3][140] , 
        \tmp[3][135] , \tmp[3][138] , \tmp[3][13] , \tmp[3][131] , 
        \tmp[3][128] , \tmp[3][11] , \tmp[3][133] , \tmp[3][137] , 
        \tmp[3][15] , n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, 
        n33, n34, n35, n36, n37, n38;
    MUX81P MX8_1_1_0 ( .D0(A[0]), .D1(A[16]), .D2(A[32]), .D3(A[48]), .D4(A
        [64]), .D5(A[80]), .D6(A[96]), .D7(A[112]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][0] ) );
    MUX81P MX8_1_1_1 ( .D0(A[1]), .D1(A[17]), .D2(A[33]), .D3(A[49]), .D4(A
        [65]), .D5(A[81]), .D6(A[97]), .D7(A[113]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][1] ) );
    MUX81P MX8_1_1_2 ( .D0(A[2]), .D1(A[18]), .D2(A[34]), .D3(A[50]), .D4(A
        [66]), .D5(A[82]), .D6(A[98]), .D7(A[114]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][2] ) );
    MUX81P MX8_1_5_10 ( .D0(A[138]), .D1(A[154]), .D2(A[170]), .D3(A[186]), 
        .D4(A[202]), .D5(A[218]), .D6(A[234]), .D7(A[250]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][138] ) );
    MUX81P MX8_1_1_3 ( .D0(A[3]), .D1(A[19]), .D2(A[35]), .D3(A[51]), .D4(A
        [67]), .D5(A[83]), .D6(A[99]), .D7(A[115]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][3] ) );
    MUX81P MX8_1_1_4 ( .D0(A[4]), .D1(A[20]), .D2(A[36]), .D3(A[52]), .D4(A
        [68]), .D5(A[84]), .D6(A[100]), .D7(A[116]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][4] ) );
    MUX81P MX8_1_1_5 ( .D0(A[5]), .D1(A[21]), .D2(A[37]), .D3(A[53]), .D4(A
        [69]), .D5(A[85]), .D6(A[101]), .D7(A[117]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][5] ) );
    MUX81P MX8_1_1_11 ( .D0(A[11]), .D1(A[27]), .D2(A[43]), .D3(A[59]), .D4(A
        [75]), .D5(A[91]), .D6(A[107]), .D7(A[123]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][11] ) );
    MUX81P MX8_1_5_3 ( .D0(A[131]), .D1(A[147]), .D2(A[163]), .D3(A[179]), 
        .D4(A[195]), .D5(A[211]), .D6(A[227]), .D7(A[243]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][131] ) );
    MUX81P MX8_1_5_4 ( .D0(A[132]), .D1(A[148]), .D2(A[164]), .D3(A[180]), 
        .D4(A[196]), .D5(A[212]), .D6(A[228]), .D7(A[244]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][132] ) );
    MUX81P MX8_1_1_10 ( .D0(A[10]), .D1(A[26]), .D2(A[42]), .D3(A[58]), .D4(A
        [74]), .D5(A[90]), .D6(A[106]), .D7(A[122]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][10] ) );
    MUX81P MX8_1_5_2 ( .D0(A[130]), .D1(A[146]), .D2(A[162]), .D3(A[178]), 
        .D4(A[194]), .D5(A[210]), .D6(A[226]), .D7(A[242]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][130] ) );
    MUX81P MX8_1_5_5 ( .D0(A[133]), .D1(A[149]), .D2(A[165]), .D3(A[181]), 
        .D4(A[197]), .D5(A[213]), .D6(A[229]), .D7(A[245]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][133] ) );
    MUX81P MX8_1_5_11 ( .D0(A[139]), .D1(A[155]), .D2(A[171]), .D3(A[187]), 
        .D4(A[203]), .D5(A[219]), .D6(A[235]), .D7(A[251]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][139] ) );
    MUX81P MX8_1_1_8 ( .D0(A[8]), .D1(A[24]), .D2(A[40]), .D3(A[56]), .D4(A
        [72]), .D5(A[88]), .D6(A[104]), .D7(A[120]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][8] ) );
    MUX81P MX8_1_5_13 ( .D0(A[141]), .D1(A[157]), .D2(A[173]), .D3(A[189]), 
        .D4(A[205]), .D5(A[221]), .D6(A[237]), .D7(A[253]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][141] ) );
    MUX81P MX8_1_1_6 ( .D0(A[6]), .D1(A[22]), .D2(A[38]), .D3(A[54]), .D4(A
        [70]), .D5(A[86]), .D6(A[102]), .D7(A[118]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][6] ) );
    MUX81P MX8_1_1_12 ( .D0(A[12]), .D1(A[28]), .D2(A[44]), .D3(A[60]), .D4(A
        [76]), .D5(A[92]), .D6(A[108]), .D7(A[124]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][12] ) );
    MUX81P MX8_1_1_15 ( .D0(A[15]), .D1(A[31]), .D2(A[47]), .D3(A[63]), .D4(A
        [79]), .D5(A[95]), .D6(A[111]), .D7(A[127]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][15] ) );
    MUX81P MX8_1_5_0 ( .D0(A[128]), .D1(A[144]), .D2(A[160]), .D3(A[176]), 
        .D4(A[192]), .D5(A[208]), .D6(A[224]), .D7(A[240]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][128] ) );
    MUX81P MX8_1_5_7 ( .D0(A[135]), .D1(A[151]), .D2(A[167]), .D3(A[183]), 
        .D4(A[199]), .D5(A[215]), .D6(A[231]), .D7(A[247]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][135] ) );
    MUX81P MX8_1_1_7 ( .D0(A[7]), .D1(A[23]), .D2(A[39]), .D3(A[55]), .D4(A
        [71]), .D5(A[87]), .D6(A[103]), .D7(A[119]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][7] ) );
    MUX81P MX8_1_5_9 ( .D0(A[137]), .D1(A[153]), .D2(A[169]), .D3(A[185]), 
        .D4(A[201]), .D5(A[217]), .D6(A[233]), .D7(A[249]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][137] ) );
    MUX81P MX8_1_5_14 ( .D0(A[142]), .D1(A[158]), .D2(A[174]), .D3(A[190]), 
        .D4(A[206]), .D5(A[222]), .D6(A[238]), .D7(A[254]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][142] ) );
    MUX81P MX8_1_1_9 ( .D0(A[9]), .D1(A[25]), .D2(A[41]), .D3(A[57]), .D4(A
        [73]), .D5(A[89]), .D6(A[105]), .D7(A[121]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][9] ) );
    MUX81P MX8_1_1_14 ( .D0(A[14]), .D1(A[30]), .D2(A[46]), .D3(A[62]), .D4(A
        [78]), .D5(A[94]), .D6(A[110]), .D7(A[126]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][14] ) );
    MUX81P MX8_1_5_1 ( .D0(A[129]), .D1(A[145]), .D2(A[161]), .D3(A[177]), 
        .D4(A[193]), .D5(A[209]), .D6(A[225]), .D7(A[241]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][129] ) );
    MUX81P MX8_1_5_8 ( .D0(A[136]), .D1(A[152]), .D2(A[168]), .D3(A[184]), 
        .D4(A[200]), .D5(A[216]), .D6(A[232]), .D7(A[248]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][136] ) );
    MUX81P MX8_1_5_15 ( .D0(A[143]), .D1(A[159]), .D2(A[175]), .D3(A[191]), 
        .D4(A[207]), .D5(A[223]), .D6(A[239]), .D7(A[255]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][143] ) );
    MUX81P MX8_1_5_12 ( .D0(A[140]), .D1(A[156]), .D2(A[172]), .D3(A[188]), 
        .D4(A[204]), .D5(A[220]), .D6(A[236]), .D7(A[252]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][140] ) );
    MUX81P MX8_1_1_13 ( .D0(A[13]), .D1(A[29]), .D2(A[45]), .D3(A[61]), .D4(A
        [77]), .D5(A[93]), .D6(A[109]), .D7(A[125]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][13] ) );
    MUX81P MX8_1_5_6 ( .D0(A[134]), .D1(A[150]), .D2(A[166]), .D3(A[182]), 
        .D4(A[198]), .D5(A[214]), .D6(A[230]), .D7(A[246]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][134] ) );
    AO2 U39 ( .A(\tmp[3][9] ), .B(n23), .C(\tmp[3][137] ), .D(SEL[3]), .Z(n22)
         );
    AO2 U40 ( .A(\tmp[3][8] ), .B(n23), .C(\tmp[3][136] ), .D(SEL[3]), .Z(n24)
         );
    AO2 U41 ( .A(\tmp[3][7] ), .B(n23), .C(\tmp[3][135] ), .D(SEL[3]), .Z(n25)
         );
    AO2 U42 ( .A(\tmp[3][6] ), .B(n23), .C(\tmp[3][134] ), .D(SEL[3]), .Z(n26)
         );
    AO2 U43 ( .A(\tmp[3][5] ), .B(n23), .C(\tmp[3][133] ), .D(SEL[3]), .Z(n27)
         );
    AO2 U44 ( .A(\tmp[3][4] ), .B(n23), .C(\tmp[3][132] ), .D(SEL[3]), .Z(n28)
         );
    AO2 U45 ( .A(\tmp[3][3] ), .B(n23), .C(\tmp[3][131] ), .D(SEL[3]), .Z(n29)
         );
    AO2 U46 ( .A(\tmp[3][2] ), .B(n23), .C(\tmp[3][130] ), .D(SEL[3]), .Z(n30)
         );
    AO2 U47 ( .A(\tmp[3][1] ), .B(n23), .C(\tmp[3][129] ), .D(SEL[3]), .Z(n31)
         );
    AO2 U48 ( .A(\tmp[3][15] ), .B(n23), .C(\tmp[3][143] ), .D(SEL[3]), .Z(n32
        ) );
    AO2 U49 ( .A(\tmp[3][14] ), .B(n23), .C(\tmp[3][142] ), .D(SEL[3]), .Z(n33
        ) );
    AO2 U50 ( .A(\tmp[3][13] ), .B(n23), .C(\tmp[3][141] ), .D(SEL[3]), .Z(n34
        ) );
    AO2 U51 ( .A(\tmp[3][12] ), .B(n23), .C(\tmp[3][140] ), .D(SEL[3]), .Z(n35
        ) );
    AO2 U52 ( .A(\tmp[3][11] ), .B(n23), .C(\tmp[3][139] ), .D(SEL[3]), .Z(n36
        ) );
    AO2 U53 ( .A(\tmp[3][10] ), .B(n23), .C(\tmp[3][138] ), .D(SEL[3]), .Z(n37
        ) );
    AO2 U54 ( .A(\tmp[3][0] ), .B(n23), .C(\tmp[3][128] ), .D(SEL[3]), .Z(n38)
         );
    IV U55 ( .A(SEL[3]), .Z(n23) );
    IV U56 ( .A(n22), .Z(MUX[9]) );
    IV U57 ( .A(n24), .Z(MUX[8]) );
    IV U58 ( .A(n25), .Z(MUX[7]) );
    IV U59 ( .A(n26), .Z(MUX[6]) );
    IV U60 ( .A(n27), .Z(MUX[5]) );
    IV U61 ( .A(n28), .Z(MUX[4]) );
    IV U62 ( .A(n29), .Z(MUX[3]) );
    IV U63 ( .A(n30), .Z(MUX[2]) );
    IV U64 ( .A(n31), .Z(MUX[1]) );
    IV U65 ( .A(n32), .Z(MUX[15]) );
    IV U66 ( .A(n33), .Z(MUX[14]) );
    IV U67 ( .A(n34), .Z(MUX[13]) );
    IV U68 ( .A(n35), .Z(MUX[12]) );
    IV U69 ( .A(n36), .Z(MUX[11]) );
    IV U70 ( .A(n37), .Z(MUX[10]) );
    IV U71 ( .A(n38), .Z(MUX[0]) );
endmodule


module fifo_DW_MEM_R_W_S_LAT_16_16_1 ( clk, wr_n, rd_addr, wr_addr, data_in, 
    data_out );
output [15:0] data_out;
input  [3:0] rd_addr;
input  [15:0] wr_addr;
input  [15:0] data_in;
input  clk, wr_n;
    wire \q[15][15] , \q[15][14] , \q[15][12] , \q[15][9] , \q[15][6] , 
        \q[15][2] , \q[14][1] , \q[10][15] , \q[6][0] , \q[1][12] , 
        \din[15][0] , \q[11][13] , \q[11][9] , \q[10][3] , \din[11][2] , 
        \din[5][1] , \din[1][3] , \q[2][2] , \din[6][12] , \q[9][14] , 
        \q[8][4] , \din[0][9] , \din[10][8] , \q[6][10] , \q[3][8] , \q[3][1] , 
        \din[10][10] , \din[8][10] , \q[0][14] , \q[11][0] , \din[10][1] , 
        \din[14][3] , \din[0][0] , \din[4][2] , \q[14][8] , \q[7][3] , 
        \din[7][14] , \din[1][10] , \q[14][5] , \q[10][7] , \q[9][10] , 
        \q[9][7] , \q[8][12] , \q[6][9] , \din[15][9] , \din[5][8] , \q[8][0] , 
        \din[10][14] , \din[8][14] , \q[2][6] , \din[11][6] , \din[0][12] , 
        \din[15][4] , \din[1][7] , \din[5][5] , \q[10][11] , \q[7][12] , 
        \q[9][3] , \q[6][4] , \din[9][12] , \q[7][7] , \din[11][12] , 
        \din[14][7] , \din[7][10] , \din[1][14] , \q[15][4] , \q[11][4] , 
        \q[8][9] , \din[10][5] , \din[4][6] , \din[0][4] , \q[7][5] , 
        \q[6][14] , \q[3][5] , \q[0][10] , \din[14][5] , \din[7][12] , 
        \din[4][4] , \q[15][0] , \q[14][7] , \q[11][15] , \q[11][6] , 
        \din[10][7] , \q[3][7] , \din[0][6] , \q[0][12] , \q[10][5] , 
        \q[9][8] , \q[9][1] , \q[8][14] , \din[11][10] , \din[9][10] , 
        \q[2][4] , \din[6][14] , \din[0][10] , \din[11][4] , \din[1][5] , 
        \din[15][6] , \q[11][11] , \q[10][13] , \q[6][6] , \din[5][7] , 
        \q[10][8] , \q[9][12] , \q[8][2] , \q[7][10] , \q[1][14] , \q[8][10] , 
        \q[2][9] , \din[11][14] , \din[9][14] , \q[9][5] , \din[1][8] , 
        \q[3][3] , \din[11][9] , \q[11][2] , \q[6][12] , \din[10][3] , 
        \din[0][2] , \din[14][1] , \q[8][6] , \q[7][1] , \din[4][0] , 
        \din[1][12] , \q[7][8] , \din[10][12] , \q[14][3] , \q[7][14] , 
        \q[1][10] , \din[14][8] , \din[8][12] , \din[4][9] , \q[6][2] , 
        \din[15][2] , \din[5][3] , \q[12][7] , \q[10][1] , \din[11][0] , 
        \q[4][4] , \q[2][0] , \din[1][1] , \wren[8] , \din[6][10] , 
        \din[0][14] , \din[5][11] , \din[3][15] , \din[7][5] , \q[0][6] , 
        \din[13][6] , \din[3][7] , \q[14][14] , \q[13][4] , \q[4][15] , 
        \q[2][11] , \q[1][5] , \din[13][13] , \din[9][1] , \din[2][13] , 
        \din[9][8] , \din[2][4] , \q[12][10] , \q[5][13] , \din[12][5] , 
        \din[6][6] , \q[14][12] , \q[14][10] , \q[13][12] , \q[13][9] , 
        \q[5][7] , \q[1][8] , \wren[1] , \din[14][11] , \din[12][15] , 
        \din[15][13] , \din[8][2] , \din[12][8] , \din[9][5] , \q[4][11] , 
        \q[2][15] , \din[2][9] , \q[12][3] , \q[0][2] , \din[3][3] , \q[4][9] , 
        \q[4][0] , \din[13][2] , \din[7][1] , \din[8][6] , \din[5][15] , 
        \din[3][11] , \wren[5] , \din[14][15] , \din[12][11] , \din[7][8] , 
        \q[13][0] , \q[12][14] , \q[5][3] , \q[3][13] , \din[6][2] , 
        \q[5][15] , \q[1][1] , \wren[13] , \din[2][0] , \din[12][1] , 
        \din[4][13] , \q[3][11] , \q[13][10] , \q[13][2] , \q[5][1] , 
        \wren[11] , \din[6][0] , \din[2][2] , \q[12][8] , \q[1][3] , 
        \din[12][3] , \din[4][11] , \din[2][15] , \din[13][9] , \q[0][9] , 
        \din[3][8] , \q[0][0] , \wren[7] , \din[12][13] , \din[8][4] , 
        \q[15][11] , \q[15][10] , \q[13][6] , \q[12][1] , \q[4][13] , 
        \q[5][8] , \q[4][2] , \din[13][0] , \din[3][1] , \din[7][3] , 
        \din[3][13] , \din[6][9] , \q[1][7] , \wren[3] , \din[15][11] , 
        \din[9][7] , \din[13][15] , \din[14][13] , \din[8][0] , \din[4][15] , 
        \din[2][11] , \q[12][12] , \wren[15] , \din[2][6] , \din[12][7] , 
        \din[6][4] , \q[12][5] , \q[5][11] , \q[3][15] , \q[5][5] , \q[4][6] , 
        \din[15][15] , \din[13][11] , \din[9][3] , \din[7][7] , \din[5][13] , 
        \din[3][5] , \q[2][13] , \din[13][4] , \q[13][15] , \q[13][14] , 
        \q[13][7] , \q[0][4] , \wren[14] , \wren[2] , \din[8][9] , 
        \din[14][12] , \din[8][1] , \q[12][13] , \q[1][6] , \din[12][6] , 
        \din[2][7] , \din[4][14] , \din[2][10] , \q[5][10] , \q[5][4] , 
        \q[3][14] , \q[4][7] , \din[15][14] , \din[6][5] , \din[13][10] , 
        \din[9][2] , \din[7][6] , \din[5][12] , \q[2][12] , \q[0][5] , 
        \din[8][8] , \q[14][13] , \q[12][4] , \din[3][4] , \q[5][14] , 
        \q[3][10] , \din[13][5] , \din[6][1] , \q[13][3] , \q[5][0] , 
        \q[1][2] , \din[4][10] , \din[2][14] , \din[2][3] , \q[12][9] , 
        \q[0][8] , \wren[10] , \din[12][2] , \din[8][5] , \din[13][8] , 
        \q[12][0] , \wren[6] , \din[12][12] , \din[3][9] , \din[13][1] , 
        \din[3][0] , \q[15][13] , \q[14][11] , \q[13][13] , \q[13][11] , 
        \q[13][8] , \q[5][9] , \q[4][12] , \q[4][3] , \q[0][1] , \din[7][2] , 
        \din[3][12] , \din[15][10] , \din[13][14] , \din[9][6] , \din[6][8] , 
        \din[12][9] , \q[12][2] , \q[1][9] , \din[15][12] , \din[2][8] , 
        \din[9][4] , \din[3][2] , \q[4][10] , \q[0][3] , \din[13][3] , 
        \q[2][14] , \q[12][15] , \q[4][8] , \q[4][1] , \din[5][14] , 
        \din[3][10] , \din[8][7] , \din[7][0] , \din[7][9] , \wren[4] , 
        \din[14][14] , \din[12][10] , \din[6][3] , \q[13][1] , \q[5][2] , 
        \q[3][12] , \q[1][0] , \din[4][12] , \wren[12] , \q[4][5] , \wren[9] , 
        \din[12][0] , \din[2][1] , \din[7][4] , \din[5][10] , \din[3][14] , 
        \q[15][8] , \q[15][1] , \q[14][15] , \q[13][5] , \q[12][6] , 
        \q[4][14] , \q[2][10] , \q[0][7] , \din[13][12] , \din[13][7] , 
        \din[3][6] , \din[9][0] , \din[2][5] , \q[5][12] , \q[1][4] , 
        \din[12][4] , \din[9][9] , \din[2][12] , \q[12][11] , \q[11][10] , 
        \q[11][3] , \q[10][9] , \q[8][11] , \q[5][6] , \din[6][7] , \wren[0] , 
        \din[14][10] , \din[12][14] , \din[8][3] , \q[9][4] , \din[9][15] , 
        \q[2][8] , \din[11][15] , \din[11][8] , \din[1][9] , \din[10][2] , 
        \din[0][3] , \q[3][2] , \q[7][0] , \q[6][13] , \din[14][0] , 
        \din[1][13] , \q[8][7] , \din[4][1] , \q[15][7] , \q[15][5] , 
        \q[14][2] , \q[7][9] , \din[14][9] , \din[8][13] , \din[4][8] , 
        \din[10][13] , \din[15][3] , \din[5][2] , \q[10][0] , \q[7][15] , 
        \q[6][3] , \q[2][1] , \q[1][11] , \din[6][11] , \din[0][15] , 
        \din[11][1] , \din[14][4] , \din[1][0] , \din[4][5] , \q[14][6] , 
        \q[11][14] , \q[7][4] , \q[3][6] , \din[7][13] , \q[0][13] , 
        \q[11][7] , \din[10][6] , \q[10][12] , \q[10][4] , \q[9][9] , 
        \q[9][0] , \din[11][11] , \din[0][7] , \q[8][15] , \din[9][11] , 
        \din[11][5] , \din[1][4] , \q[2][5] , \din[6][15] , \din[0][11] , 
        \q[7][11] , \q[1][15] , \q[6][7] , \din[15][7] , \q[14][4] , 
        \q[10][10] , \q[10][6] , \q[9][13] , \q[8][3] , \din[5][6] , 
        \q[9][11] , \q[8][1] , \din[10][15] , \din[8][15] , \din[11][7] , 
        \q[7][13] , \q[6][5] , \q[2][7] , \din[1][6] , \din[0][13] , 
        \din[15][5] , \din[5][4] , \q[9][2] , \din[11][13] , \din[9][13] , 
        \din[14][6] , \q[15][3] , \q[14][0] , \q[11][5] , \q[8][8] , \q[7][6] , 
        \din[4][7] , \q[6][15] , \q[3][4] , \din[7][11] , \din[1][15] , 
        \q[0][11] , \din[10][4] , \din[0][5] , \din[15][1] , \q[11][12] , 
        \q[11][8] , \q[10][14] , \din[5][0] , \q[10][2] , \q[6][1] , 
        \q[1][13] , \q[2][3] , \din[11][3] , \din[6][13] , \din[1][2] , 
        \q[3][9] , \q[11][1] , \q[9][15] , \q[8][5] , \din[0][8] , 
        \din[10][11] , \din[10][9] , \din[8][11] , \din[10][0] , \q[6][11] , 
        \q[3][0] , \din[0][1] , \q[0][15] , \q[7][2] , \din[14][2] , 
        \din[7][15] , \din[1][11] , \din[4][3] , \q[14][9] , \q[6][8] , 
        \q[9][6] , \q[8][13] , \din[15][8] , \din[5][9] , n38, n39, n40, n41, 
        n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54;
    fifo_DW01_mux_any_256_4_16_1 MX ( .A({\q[15][15] , \q[15][14] , 
        \q[15][13] , \q[15][12] , \q[15][11] , \q[15][10] , \q[15][9] , 
        \q[15][8] , \q[15][7] , \q[15][6] , \q[15][5] , \q[15][4] , \q[15][3] , 
        \q[15][2] , \q[15][1] , \q[15][0] , \q[14][15] , \q[14][14] , 
        \q[14][13] , \q[14][12] , \q[14][11] , \q[14][10] , \q[14][9] , 
        \q[14][8] , \q[14][7] , \q[14][6] , \q[14][5] , \q[14][4] , \q[14][3] , 
        \q[14][2] , \q[14][1] , \q[14][0] , \q[13][15] , \q[13][14] , 
        \q[13][13] , \q[13][12] , \q[13][11] , \q[13][10] , \q[13][9] , 
        \q[13][8] , \q[13][7] , \q[13][6] , \q[13][5] , \q[13][4] , \q[13][3] , 
        \q[13][2] , \q[13][1] , \q[13][0] , \q[12][15] , \q[12][14] , 
        \q[12][13] , \q[12][12] , \q[12][11] , \q[12][10] , \q[12][9] , 
        \q[12][8] , \q[12][7] , \q[12][6] , \q[12][5] , \q[12][4] , \q[12][3] , 
        \q[12][2] , \q[12][1] , \q[12][0] , \q[11][15] , \q[11][14] , 
        \q[11][13] , \q[11][12] , \q[11][11] , \q[11][10] , \q[11][9] , 
        \q[11][8] , \q[11][7] , \q[11][6] , \q[11][5] , \q[11][4] , \q[11][3] , 
        \q[11][2] , \q[11][1] , \q[11][0] , \q[10][15] , \q[10][14] , 
        \q[10][13] , \q[10][12] , \q[10][11] , \q[10][10] , \q[10][9] , 
        \q[10][8] , \q[10][7] , \q[10][6] , \q[10][5] , \q[10][4] , \q[10][3] , 
        \q[10][2] , \q[10][1] , \q[10][0] , \q[9][15] , \q[9][14] , \q[9][13] , 
        \q[9][12] , \q[9][11] , \q[9][10] , \q[9][9] , \q[9][8] , \q[9][7] , 
        \q[9][6] , \q[9][5] , \q[9][4] , \q[9][3] , \q[9][2] , \q[9][1] , 
        \q[9][0] , \q[8][15] , \q[8][14] , \q[8][13] , \q[8][12] , \q[8][11] , 
        \q[8][10] , \q[8][9] , \q[8][8] , \q[8][7] , \q[8][6] , \q[8][5] , 
        \q[8][4] , \q[8][3] , \q[8][2] , \q[8][1] , \q[8][0] , \q[7][15] , 
        \q[7][14] , \q[7][13] , \q[7][12] , \q[7][11] , \q[7][10] , \q[7][9] , 
        \q[7][8] , \q[7][7] , \q[7][6] , \q[7][5] , \q[7][4] , \q[7][3] , 
        \q[7][2] , \q[7][1] , \q[7][0] , \q[6][15] , \q[6][14] , \q[6][13] , 
        \q[6][12] , \q[6][11] , \q[6][10] , \q[6][9] , \q[6][8] , \q[6][7] , 
        \q[6][6] , \q[6][5] , \q[6][4] , \q[6][3] , \q[6][2] , \q[6][1] , 
        \q[6][0] , \q[5][15] , \q[5][14] , \q[5][13] , \q[5][12] , \q[5][11] , 
        \q[5][10] , \q[5][9] , \q[5][8] , \q[5][7] , \q[5][6] , \q[5][5] , 
        \q[5][4] , \q[5][3] , \q[5][2] , \q[5][1] , \q[5][0] , \q[4][15] , 
        \q[4][14] , \q[4][13] , \q[4][12] , \q[4][11] , \q[4][10] , \q[4][9] , 
        \q[4][8] , \q[4][7] , \q[4][6] , \q[4][5] , \q[4][4] , \q[4][3] , 
        \q[4][2] , \q[4][1] , \q[4][0] , \q[3][15] , \q[3][14] , \q[3][13] , 
        \q[3][12] , \q[3][11] , \q[3][10] , \q[3][9] , \q[3][8] , \q[3][7] , 
        \q[3][6] , \q[3][5] , \q[3][4] , \q[3][3] , \q[3][2] , \q[3][1] , 
        \q[3][0] , \q[2][15] , \q[2][14] , \q[2][13] , \q[2][12] , \q[2][11] , 
        \q[2][10] , \q[2][9] , \q[2][8] , \q[2][7] , \q[2][6] , \q[2][5] , 
        \q[2][4] , \q[2][3] , \q[2][2] , \q[2][1] , \q[2][0] , \q[1][15] , 
        \q[1][14] , \q[1][13] , \q[1][12] , \q[1][11] , \q[1][10] , \q[1][9] , 
        \q[1][8] , \q[1][7] , \q[1][6] , \q[1][5] , \q[1][4] , \q[1][3] , 
        \q[1][2] , \q[1][1] , \q[1][0] , \q[0][15] , \q[0][14] , \q[0][13] , 
        \q[0][12] , \q[0][11] , \q[0][10] , \q[0][9] , \q[0][8] , \q[0][7] , 
        \q[0][6] , \q[0][5] , \q[0][4] , \q[0][3] , \q[0][2] , \q[0][1] , 
        \q[0][0] }), .SEL(rd_addr), .MUX(data_out) );
    MUX21H MX1_0_0 ( .A(\q[0][0] ), .B(data_in[0]), .S(\wren[0] ), .Z(
        \din[0][0] ) );
    MUX21H MX1_0_11 ( .A(\q[11][0] ), .B(data_in[0]), .S(\wren[11] ), .Z(
        \din[11][0] ) );
    MUX21H MX1_8_1 ( .A(\q[1][8] ), .B(data_in[8]), .S(\wren[1] ), .Z(
        \din[1][8] ) );
    MUX21H MX1_15_9 ( .A(\q[9][15] ), .B(data_in[15]), .S(\wren[9] ), .Z(
        \din[9][15] ) );
    MUX21H MX1_12_3 ( .A(\q[3][12] ), .B(data_in[12]), .S(\wren[3] ), .Z(
        \din[3][12] ) );
    MUX21H MX1_14_12 ( .A(\q[12][14] ), .B(data_in[14]), .S(\wren[12] ), .Z(
        \din[12][14] ) );
    MUX21H MX1_5_6 ( .A(\q[6][5] ), .B(data_in[5]), .S(\wren[6] ), .Z(
        \din[6][5] ) );
    MUX21H MX1_6_14 ( .A(\q[14][6] ), .B(data_in[6]), .S(\wren[14] ), .Z(
        \din[14][6] ) );
    MUX21H MX1_1_0 ( .A(\q[0][1] ), .B(data_in[1]), .S(\wren[0] ), .Z(
        \din[0][1] ) );
    MUX21H MX1_4_6 ( .A(\q[6][4] ), .B(data_in[4]), .S(\wren[6] ), .Z(
        \din[6][4] ) );
    MUX21H MX1_1_10 ( .A(\q[10][1] ), .B(data_in[1]), .S(\wren[10] ), .Z(
        \din[10][1] ) );
    MUX21H MX1_0_9 ( .A(\q[9][0] ), .B(data_in[0]), .S(\wren[9] ), .Z(
        \din[9][0] ) );
    MUX21H MX1_4_10 ( .A(\q[10][4] ), .B(data_in[4]), .S(\wren[10] ), .Z(
        \din[10][4] ) );
    MUX21H MX1_14_9 ( .A(\q[9][14] ), .B(data_in[14]), .S(\wren[9] ), .Z(
        \din[9][14] ) );
    MUX21H MX1_7_15 ( .A(\q[15][7] ), .B(data_in[7]), .S(\wren[15] ), .Z(
        \din[15][7] ) );
    MUX21H MX1_15_13 ( .A(\q[13][15] ), .B(data_in[15]), .S(\wren[13] ), .Z(
        \din[13][15] ) );
    MUX21H MX1_9_1 ( .A(\q[1][9] ), .B(data_in[9]), .S(\wren[1] ), .Z(
        \din[1][9] ) );
    MUX21H MX1_8_8 ( .A(\q[8][8] ), .B(data_in[8]), .S(\wren[8] ), .Z(
        \din[8][8] ) );
    MUX21H MX1_13_3 ( .A(\q[3][13] ), .B(data_in[13]), .S(\wren[3] ), .Z(
        \din[3][13] ) );
    MUX21H MX1_15_0 ( .A(\q[0][15] ), .B(data_in[15]), .S(\wren[0] ), .Z(
        \din[0][15] ) );
    MUX21H MX1_10_6 ( .A(\q[6][10] ), .B(data_in[10]), .S(\wren[6] ), .Z(
        \din[6][10] ) );
    MUX21H MX1_1_9 ( .A(\q[9][1] ), .B(data_in[1]), .S(\wren[9] ), .Z(
        \din[9][1] ) );
    MUX21H MX1_2_5 ( .A(\q[5][2] ), .B(data_in[2]), .S(\wren[5] ), .Z(
        \din[5][2] ) );
    MUX21H MX1_8_13 ( .A(\q[13][8] ), .B(data_in[8]), .S(\wren[13] ), .Z(
        \din[13][8] ) );
    MUX21H MX1_2_15 ( .A(\q[15][2] ), .B(data_in[2]), .S(\wren[15] ), .Z(
        \din[15][2] ) );
    MUX21H MX1_7_3 ( .A(\q[3][7] ), .B(data_in[7]), .S(\wren[3] ), .Z(
        \din[3][7] ) );
    MUX21H MX1_10_13 ( .A(\q[13][10] ), .B(data_in[10]), .S(\wren[13] ), .Z(
        \din[13][10] ) );
    MUX21H MX1_5_11 ( .A(\q[11][5] ), .B(data_in[5]), .S(\wren[11] ), .Z(
        \din[11][5] ) );
    MUX21H MX1_6_3 ( .A(\q[3][6] ), .B(data_in[6]), .S(\wren[3] ), .Z(
        \din[3][6] ) );
    MUX21H MX1_3_5 ( .A(\q[5][3] ), .B(data_in[3]), .S(\wren[5] ), .Z(
        \din[5][3] ) );
    MUX21H MX1_3_14 ( .A(\q[14][3] ), .B(data_in[3]), .S(\wren[14] ), .Z(
        \din[14][3] ) );
    MUX21H MX1_9_8 ( .A(\q[8][9] ), .B(data_in[9]), .S(\wren[8] ), .Z(
        \din[8][9] ) );
    MUX21H MX1_9_12 ( .A(\q[12][9] ), .B(data_in[9]), .S(\wren[12] ), .Z(
        \din[12][9] ) );
    MUX21H MX1_11_6 ( .A(\q[6][11] ), .B(data_in[11]), .S(\wren[6] ), .Z(
        \din[6][11] ) );
    MUX21H MX1_14_0 ( .A(\q[0][14] ), .B(data_in[14]), .S(\wren[0] ), .Z(
        \din[0][14] ) );
    MUX21H MX1_9_15 ( .A(\q[15][9] ), .B(data_in[9]), .S(\wren[15] ), .Z(
        \din[15][9] ) );
    MUX21H MX1_11_12 ( .A(\q[12][11] ), .B(data_in[11]), .S(\wren[12] ), .Z(
        \din[12][11] ) );
    MUX21H MX1_14_7 ( .A(\q[7][14] ), .B(data_in[14]), .S(\wren[7] ), .Z(
        \din[7][14] ) );
    MUX21H MX1_11_1 ( .A(\q[1][11] ), .B(data_in[11]), .S(\wren[1] ), .Z(
        \din[1][11] ) );
    MUX21H MX1_3_13 ( .A(\q[13][3] ), .B(data_in[3]), .S(\wren[13] ), .Z(
        \din[13][3] ) );
    MUX21H MX1_11_15 ( .A(\q[15][11] ), .B(data_in[11]), .S(\wren[15] ), .Z(
        \din[15][11] ) );
    MUX21H MX1_4_8 ( .A(\q[8][4] ), .B(data_in[4]), .S(\wren[8] ), .Z(
        \din[8][4] ) );
    MUX21H MX1_3_2 ( .A(\q[2][3] ), .B(data_in[3]), .S(\wren[2] ), .Z(
        \din[2][3] ) );
    MUX21H MX1_6_4 ( .A(\q[4][6] ), .B(data_in[6]), .S(\wren[4] ), .Z(
        \din[4][6] ) );
    MUX21H MX1_2_2 ( .A(\q[2][2] ), .B(data_in[2]), .S(\wren[2] ), .Z(
        \din[2][2] ) );
    MUX21H MX1_2_12 ( .A(\q[12][2] ), .B(data_in[2]), .S(\wren[12] ), .Z(
        \din[12][2] ) );
    MUX21H MX1_5_8 ( .A(\q[8][5] ), .B(data_in[5]), .S(\wren[8] ), .Z(
        \din[8][5] ) );
    MUX21H MX1_8_14 ( .A(\q[14][8] ), .B(data_in[8]), .S(\wren[14] ), .Z(
        \din[14][8] ) );
    MUX21H MX1_10_14 ( .A(\q[14][10] ), .B(data_in[10]), .S(\wren[14] ), .Z(
        \din[14][10] ) );
    MUX21H MX1_7_4 ( .A(\q[4][7] ), .B(data_in[7]), .S(\wren[4] ), .Z(
        \din[4][7] ) );
    MUX21H MX1_7_12 ( .A(\q[12][7] ), .B(data_in[7]), .S(\wren[12] ), .Z(
        \din[12][7] ) );
    MUX21H MX1_10_1 ( .A(\q[1][10] ), .B(data_in[10]), .S(\wren[1] ), .Z(
        \din[1][10] ) );
    MUX21H MX1_15_7 ( .A(\q[7][15] ), .B(data_in[15]), .S(\wren[7] ), .Z(
        \din[7][15] ) );
    MUX21H MX1_9_6 ( .A(\q[6][9] ), .B(data_in[9]), .S(\wren[6] ), .Z(
        \din[6][9] ) );
    MUX21H MX1_11_8 ( .A(\q[8][11] ), .B(data_in[11]), .S(\wren[8] ), .Z(
        \din[8][11] ) );
    MUX21H MX1_13_4 ( .A(\q[4][13] ), .B(data_in[13]), .S(\wren[4] ), .Z(
        \din[4][13] ) );
    MUX21H MX1_15_14 ( .A(\q[14][15] ), .B(data_in[15]), .S(\wren[14] ), .Z(
        \din[14][15] ) );
    MUX21H MX1_0_1 ( .A(\q[1][0] ), .B(data_in[0]), .S(\wren[1] ), .Z(
        \din[1][0] ) );
    MUX21H MX1_0_6 ( .A(\q[6][0] ), .B(data_in[0]), .S(\wren[6] ), .Z(
        \din[6][0] ) );
    MUX21H MX1_0_7 ( .A(\q[7][0] ), .B(data_in[0]), .S(\wren[7] ), .Z(
        \din[7][0] ) );
    MUX21H MX1_1_7 ( .A(\q[7][1] ), .B(data_in[1]), .S(\wren[7] ), .Z(
        \din[7][1] ) );
    MUX21H MX1_4_1 ( .A(\q[1][4] ), .B(data_in[4]), .S(\wren[1] ), .Z(
        \din[1][4] ) );
    MUX21H MX1_13_11 ( .A(\q[11][13] ), .B(data_in[13]), .S(\wren[11] ), .Z(
        \din[11][13] ) );
    MUX21H MX1_5_1 ( .A(\q[1][5] ), .B(data_in[5]), .S(\wren[1] ), .Z(
        \din[1][5] ) );
    MUX21H MX1_6_13 ( .A(\q[13][6] ), .B(data_in[6]), .S(\wren[13] ), .Z(
        \din[13][6] ) );
    MUX21H MX1_14_15 ( .A(\q[15][14] ), .B(data_in[14]), .S(\wren[15] ), .Z(
        \din[15][14] ) );
    MUX21H MX1_8_6 ( .A(\q[6][8] ), .B(data_in[8]), .S(\wren[6] ), .Z(
        \din[6][8] ) );
    MUX21H MX1_8_15 ( .A(\q[15][8] ), .B(data_in[8]), .S(\wren[15] ), .Z(
        \din[15][8] ) );
    MUX21H MX1_10_8 ( .A(\q[8][10] ), .B(data_in[10]), .S(\wren[8] ), .Z(
        \din[8][10] ) );
    MUX21H MX1_12_10 ( .A(\q[10][12] ), .B(data_in[12]), .S(\wren[10] ), .Z(
        \din[10][12] ) );
    MUX21H MX1_12_4 ( .A(\q[4][12] ), .B(data_in[12]), .S(\wren[4] ), .Z(
        \din[4][12] ) );
    MUX21H MX1_10_0 ( .A(\q[0][10] ), .B(data_in[10]), .S(\wren[0] ), .Z(
        \din[0][10] ) );
    MUX21H MX1_15_6 ( .A(\q[6][15] ), .B(data_in[15]), .S(\wren[6] ), .Z(
        \din[6][15] ) );
    MUX21H MX1_2_3 ( .A(\q[3][2] ), .B(data_in[2]), .S(\wren[3] ), .Z(
        \din[3][2] ) );
    MUX21H MX1_2_13 ( .A(\q[13][2] ), .B(data_in[2]), .S(\wren[13] ), .Z(
        \din[13][2] ) );
    MUX21H MX1_5_9 ( .A(\q[9][5] ), .B(data_in[5]), .S(\wren[9] ), .Z(
        \din[9][5] ) );
    MUX21H MX1_7_5 ( .A(\q[5][7] ), .B(data_in[7]), .S(\wren[5] ), .Z(
        \din[5][7] ) );
    MUX21H MX1_10_15 ( .A(\q[15][10] ), .B(data_in[10]), .S(\wren[15] ), .Z(
        \din[15][10] ) );
    MUX21H MX1_4_9 ( .A(\q[9][4] ), .B(data_in[4]), .S(\wren[9] ), .Z(
        \din[9][4] ) );
    MUX21H MX1_3_3 ( .A(\q[3][3] ), .B(data_in[3]), .S(\wren[3] ), .Z(
        \din[3][3] ) );
    MUX21H MX1_6_5 ( .A(\q[5][6] ), .B(data_in[6]), .S(\wren[5] ), .Z(
        \din[5][6] ) );
    MUX21H MX1_9_14 ( .A(\q[14][9] ), .B(data_in[9]), .S(\wren[14] ), .Z(
        \din[14][9] ) );
    MUX21H MX1_14_6 ( .A(\q[6][14] ), .B(data_in[14]), .S(\wren[6] ), .Z(
        \din[6][14] ) );
    MUX21H MX1_11_0 ( .A(\q[0][11] ), .B(data_in[11]), .S(\wren[0] ), .Z(
        \din[0][11] ) );
    MUX21H MX1_3_12 ( .A(\q[12][3] ), .B(data_in[3]), .S(\wren[12] ), .Z(
        \din[12][3] ) );
    MUX21H MX1_11_14 ( .A(\q[14][11] ), .B(data_in[11]), .S(\wren[14] ), .Z(
        \din[14][11] ) );
    MUX21H MX1_5_0 ( .A(\q[0][5] ), .B(data_in[5]), .S(\wren[0] ), .Z(
        \din[0][5] ) );
    MUX21H MX1_8_7 ( .A(\q[7][8] ), .B(data_in[8]), .S(\wren[7] ), .Z(
        \din[7][8] ) );
    MUX21H MX1_10_9 ( .A(\q[9][10] ), .B(data_in[10]), .S(\wren[9] ), .Z(
        \din[9][10] ) );
    MUX21H MX1_12_11 ( .A(\q[11][12] ), .B(data_in[12]), .S(\wren[11] ), .Z(
        \din[11][12] ) );
    MUX21H MX1_12_5 ( .A(\q[5][12] ), .B(data_in[12]), .S(\wren[5] ), .Z(
        \din[5][12] ) );
    MUX21H MX1_6_12 ( .A(\q[12][6] ), .B(data_in[6]), .S(\wren[12] ), .Z(
        \din[12][6] ) );
    MUX21H MX1_14_14 ( .A(\q[14][14] ), .B(data_in[14]), .S(\wren[14] ), .Z(
        \din[14][14] ) );
    MUX21H MX1_1_6 ( .A(\q[6][1] ), .B(data_in[1]), .S(\wren[6] ), .Z(
        \din[6][1] ) );
    MUX21H MX1_4_0 ( .A(\q[0][4] ), .B(data_in[4]), .S(\wren[0] ), .Z(
        \din[0][4] ) );
    MUX21H MX1_7_13 ( .A(\q[13][7] ), .B(data_in[7]), .S(\wren[13] ), .Z(
        \din[13][7] ) );
    MUX21H MX1_13_10 ( .A(\q[10][13] ), .B(data_in[13]), .S(\wren[10] ), .Z(
        \din[10][13] ) );
    MUX21H MX1_11_9 ( .A(\q[9][11] ), .B(data_in[11]), .S(\wren[9] ), .Z(
        \din[9][11] ) );
    MUX21H MX1_9_7 ( .A(\q[7][9] ), .B(data_in[9]), .S(\wren[7] ), .Z(
        \din[7][9] ) );
    MUX21H MX1_13_5 ( .A(\q[5][13] ), .B(data_in[13]), .S(\wren[5] ), .Z(
        \din[5][13] ) );
    MUX21H MX1_15_15 ( .A(\q[15][15] ), .B(data_in[15]), .S(\wren[15] ), .Z(
        \din[15][15] ) );
    MUX21H MX1_7_14 ( .A(\q[14][7] ), .B(data_in[7]), .S(\wren[14] ), .Z(
        \din[14][7] ) );
    MUX21H MX1_9_0 ( .A(\q[0][9] ), .B(data_in[9]), .S(\wren[0] ), .Z(
        \din[0][9] ) );
    MUX21H MX1_14_8 ( .A(\q[8][14] ), .B(data_in[14]), .S(\wren[8] ), .Z(
        \din[8][14] ) );
    MUX21H MX1_15_12 ( .A(\q[12][15] ), .B(data_in[15]), .S(\wren[12] ), .Z(
        \din[12][15] ) );
    MUX21H MX1_13_2 ( .A(\q[2][13] ), .B(data_in[13]), .S(\wren[2] ), .Z(
        \din[2][13] ) );
    MUX21H MX1_1_1 ( .A(\q[1][1] ), .B(data_in[1]), .S(\wren[1] ), .Z(
        \din[1][1] ) );
    MUX21H MX1_1_11 ( .A(\q[11][1] ), .B(data_in[1]), .S(\wren[11] ), .Z(
        \din[11][1] ) );
    MUX21H MX1_4_7 ( .A(\q[7][4] ), .B(data_in[4]), .S(\wren[7] ), .Z(
        \din[7][4] ) );
    MUX21H MX1_14_13 ( .A(\q[13][14] ), .B(data_in[14]), .S(\wren[13] ), .Z(
        \din[13][14] ) );
    MUX21H MX1_0_2 ( .A(\q[2][0] ), .B(data_in[0]), .S(\wren[2] ), .Z(
        \din[2][0] ) );
    MUX21H MX1_0_3 ( .A(\q[3][0] ), .B(data_in[0]), .S(\wren[3] ), .Z(
        \din[3][0] ) );
    MUX21H MX1_0_8 ( .A(\q[8][0] ), .B(data_in[0]), .S(\wren[8] ), .Z(
        \din[8][0] ) );
    MUX21H MX1_0_10 ( .A(\q[10][0] ), .B(data_in[0]), .S(\wren[10] ), .Z(
        \din[10][0] ) );
    MUX21H MX1_5_7 ( .A(\q[7][5] ), .B(data_in[5]), .S(\wren[7] ), .Z(
        \din[7][5] ) );
    MUX21H MX1_6_15 ( .A(\q[15][6] ), .B(data_in[6]), .S(\wren[15] ), .Z(
        \din[15][6] ) );
    MUX21H MX1_8_0 ( .A(\q[0][8] ), .B(data_in[8]), .S(\wren[0] ), .Z(
        \din[0][8] ) );
    MUX21H MX1_1_8 ( .A(\q[8][1] ), .B(data_in[1]), .S(\wren[8] ), .Z(
        \din[8][1] ) );
    MUX21H MX1_3_15 ( .A(\q[15][3] ), .B(data_in[3]), .S(\wren[15] ), .Z(
        \din[15][3] ) );
    MUX21H MX1_12_2 ( .A(\q[2][12] ), .B(data_in[12]), .S(\wren[2] ), .Z(
        \din[2][12] ) );
    MUX21H MX1_15_8 ( .A(\q[8][15] ), .B(data_in[15]), .S(\wren[8] ), .Z(
        \din[8][15] ) );
    MUX21H MX1_9_9 ( .A(\q[9][9] ), .B(data_in[9]), .S(\wren[9] ), .Z(
        \din[9][9] ) );
    MUX21H MX1_11_7 ( .A(\q[7][11] ), .B(data_in[11]), .S(\wren[7] ), .Z(
        \din[7][11] ) );
    MUX21H MX1_9_13 ( .A(\q[13][9] ), .B(data_in[9]), .S(\wren[13] ), .Z(
        \din[13][9] ) );
    MUX21H MX1_14_1 ( .A(\q[1][14] ), .B(data_in[14]), .S(\wren[1] ), .Z(
        \din[1][14] ) );
    MUX21H MX1_11_13 ( .A(\q[13][11] ), .B(data_in[11]), .S(\wren[13] ), .Z(
        \din[13][11] ) );
    MUX21H MX1_5_10 ( .A(\q[10][5] ), .B(data_in[5]), .S(\wren[10] ), .Z(
        \din[10][5] ) );
    MUX21H MX1_6_2 ( .A(\q[2][6] ), .B(data_in[6]), .S(\wren[2] ), .Z(
        \din[2][6] ) );
    MUX21H MX1_3_4 ( .A(\q[4][3] ), .B(data_in[3]), .S(\wren[4] ), .Z(
        \din[4][3] ) );
    MUX21H MX1_0_12 ( .A(\q[12][0] ), .B(data_in[0]), .S(\wren[12] ), .Z(
        \din[12][0] ) );
    MUX21H MX1_2_4 ( .A(\q[4][2] ), .B(data_in[2]), .S(\wren[4] ), .Z(
        \din[4][2] ) );
    MUX21H MX1_8_12 ( .A(\q[12][8] ), .B(data_in[8]), .S(\wren[12] ), .Z(
        \din[12][8] ) );
    MUX21H MX1_2_14 ( .A(\q[14][2] ), .B(data_in[2]), .S(\wren[14] ), .Z(
        \din[14][2] ) );
    MUX21H MX1_7_2 ( .A(\q[2][7] ), .B(data_in[7]), .S(\wren[2] ), .Z(
        \din[2][7] ) );
    MUX21H MX1_4_11 ( .A(\q[11][4] ), .B(data_in[4]), .S(\wren[11] ), .Z(
        \din[11][4] ) );
    MUX21H MX1_10_12 ( .A(\q[12][10] ), .B(data_in[10]), .S(\wren[12] ), .Z(
        \din[12][10] ) );
    MUX21H MX1_8_9 ( .A(\q[9][8] ), .B(data_in[8]), .S(\wren[9] ), .Z(
        \din[9][8] ) );
    MUX21H MX1_10_7 ( .A(\q[7][10] ), .B(data_in[10]), .S(\wren[7] ), .Z(
        \din[7][10] ) );
    MUX21H MX1_15_1 ( .A(\q[1][15] ), .B(data_in[15]), .S(\wren[1] ), .Z(
        \din[1][15] ) );
    MUX21H MX1_12_0 ( .A(\q[0][12] ), .B(data_in[12]), .S(\wren[0] ), .Z(
        \din[0][12] ) );
    MUX21H MX1_8_2 ( .A(\q[2][8] ), .B(data_in[8]), .S(\wren[2] ), .Z(
        \din[2][8] ) );
    MUX21H MX1_12_14 ( .A(\q[14][12] ), .B(data_in[12]), .S(\wren[14] ), .Z(
        \din[14][12] ) );
    MUX21H MX1_7_9 ( .A(\q[9][7] ), .B(data_in[7]), .S(\wren[9] ), .Z(
        \din[9][7] ) );
    MUX21H MX1_5_5 ( .A(\q[5][5] ), .B(data_in[5]), .S(\wren[5] ), .Z(
        \din[5][5] ) );
    MUX21H MX1_1_3 ( .A(\q[3][1] ), .B(data_in[1]), .S(\wren[3] ), .Z(
        \din[3][1] ) );
    MUX21H MX1_6_9 ( .A(\q[9][6] ), .B(data_in[6]), .S(\wren[9] ), .Z(
        \din[9][6] ) );
    MUX21H MX1_14_11 ( .A(\q[11][14] ), .B(data_in[14]), .S(\wren[11] ), .Z(
        \din[11][14] ) );
    MUX21H MX1_1_13 ( .A(\q[13][1] ), .B(data_in[1]), .S(\wren[13] ), .Z(
        \din[13][1] ) );
    MUX21H MX1_2_1 ( .A(\q[1][2] ), .B(data_in[2]), .S(\wren[1] ), .Z(
        \din[1][2] ) );
    MUX21H MX1_2_6 ( .A(\q[6][2] ), .B(data_in[2]), .S(\wren[6] ), .Z(
        \din[6][2] ) );
    MUX21H MX1_4_5 ( .A(\q[5][4] ), .B(data_in[4]), .S(\wren[5] ), .Z(
        \din[5][4] ) );
    MUX21H MX1_13_15 ( .A(\q[15][13] ), .B(data_in[13]), .S(\wren[15] ), .Z(
        \din[15][13] ) );
    MUX21H MX1_4_13 ( .A(\q[13][4] ), .B(data_in[4]), .S(\wren[13] ), .Z(
        \din[13][4] ) );
    MUX21H MX1_9_2 ( .A(\q[2][9] ), .B(data_in[9]), .S(\wren[2] ), .Z(
        \din[2][9] ) );
    MUX21H MX1_13_0 ( .A(\q[0][13] ), .B(data_in[13]), .S(\wren[0] ), .Z(
        \din[0][13] ) );
    MUX21H MX1_15_10 ( .A(\q[10][15] ), .B(data_in[15]), .S(\wren[10] ), .Z(
        \din[10][15] ) );
    MUX21H MX1_12_9 ( .A(\q[9][12] ), .B(data_in[12]), .S(\wren[9] ), .Z(
        \din[9][12] ) );
    MUX21H MX1_7_0 ( .A(\q[0][7] ), .B(data_in[7]), .S(\wren[0] ), .Z(
        \din[0][7] ) );
    MUX21H MX1_10_5 ( .A(\q[5][10] ), .B(data_in[10]), .S(\wren[5] ), .Z(
        \din[5][10] ) );
    MUX21H MX1_15_3 ( .A(\q[3][15] ), .B(data_in[15]), .S(\wren[3] ), .Z(
        \din[3][15] ) );
    MUX21H MX1_10_10 ( .A(\q[10][10] ), .B(data_in[10]), .S(\wren[10] ), .Z(
        \din[10][10] ) );
    MUX21H MX1_8_10 ( .A(\q[10][8] ), .B(data_in[8]), .S(\wren[10] ), .Z(
        \din[10][8] ) );
    MUX21H MX1_3_6 ( .A(\q[6][3] ), .B(data_in[3]), .S(\wren[6] ), .Z(
        \din[6][3] ) );
    MUX21H MX1_3_10 ( .A(\q[10][3] ), .B(data_in[3]), .S(\wren[10] ), .Z(
        \din[10][3] ) );
    MUX21H MX1_5_12 ( .A(\q[12][5] ), .B(data_in[5]), .S(\wren[12] ), .Z(
        \din[12][5] ) );
    MUX21H MX1_6_0 ( .A(\q[0][6] ), .B(data_in[6]), .S(\wren[0] ), .Z(
        \din[0][6] ) );
    MUX21H MX1_9_11 ( .A(\q[11][9] ), .B(data_in[9]), .S(\wren[11] ), .Z(
        \din[11][9] ) );
    MUX21H MX1_11_11 ( .A(\q[11][11] ), .B(data_in[11]), .S(\wren[11] ), .Z(
        \din[11][11] ) );
    MUX21H MX1_13_9 ( .A(\q[9][13] ), .B(data_in[13]), .S(\wren[9] ), .Z(
        \din[9][13] ) );
    MUX21H MX1_14_3 ( .A(\q[3][14] ), .B(data_in[14]), .S(\wren[3] ), .Z(
        \din[3][14] ) );
    MUX21H MX1_11_5 ( .A(\q[5][11] ), .B(data_in[11]), .S(\wren[5] ), .Z(
        \din[5][11] ) );
    MUX21H MX1_3_1 ( .A(\q[1][3] ), .B(data_in[3]), .S(\wren[1] ), .Z(
        \din[1][3] ) );
    MUX21H MX1_5_15 ( .A(\q[15][5] ), .B(data_in[5]), .S(\wren[15] ), .Z(
        \din[15][5] ) );
    MUX21H MX1_6_7 ( .A(\q[7][6] ), .B(data_in[6]), .S(\wren[7] ), .Z(
        \din[7][6] ) );
    MUX21H MX1_11_2 ( .A(\q[2][11] ), .B(data_in[11]), .S(\wren[2] ), .Z(
        \din[2][11] ) );
    MUX21H MX1_14_4 ( .A(\q[4][14] ), .B(data_in[14]), .S(\wren[4] ), .Z(
        \din[4][14] ) );
    MUX21H MX1_2_11 ( .A(\q[11][2] ), .B(data_in[2]), .S(\wren[11] ), .Z(
        \din[11][2] ) );
    MUX21H MX1_3_8 ( .A(\q[8][3] ), .B(data_in[3]), .S(\wren[8] ), .Z(
        \din[8][3] ) );
    MUX21H MX1_4_14 ( .A(\q[14][4] ), .B(data_in[4]), .S(\wren[14] ), .Z(
        \din[14][4] ) );
    MUX21H MX1_7_7 ( .A(\q[7][7] ), .B(data_in[7]), .S(\wren[7] ), .Z(
        \din[7][7] ) );
    MUX21H MX1_10_2 ( .A(\q[2][10] ), .B(data_in[10]), .S(\wren[2] ), .Z(
        \din[2][10] ) );
    MUX21H MX1_15_4 ( .A(\q[4][15] ), .B(data_in[15]), .S(\wren[4] ), .Z(
        \din[4][15] ) );
    MUX21H MX1_13_7 ( .A(\q[7][13] ), .B(data_in[13]), .S(\wren[7] ), .Z(
        \din[7][13] ) );
    MUX21H MX1_7_11 ( .A(\q[11][7] ), .B(data_in[7]), .S(\wren[11] ), .Z(
        \din[11][7] ) );
    MUX21H MX1_9_5 ( .A(\q[5][9] ), .B(data_in[9]), .S(\wren[5] ), .Z(
        \din[5][9] ) );
    MUX21H MX1_4_2 ( .A(\q[2][4] ), .B(data_in[4]), .S(\wren[2] ), .Z(
        \din[2][4] ) );
    MUX21H MX1_13_12 ( .A(\q[12][13] ), .B(data_in[13]), .S(\wren[12] ), .Z(
        \din[12][13] ) );
    MUX21H MX1_0_4 ( .A(\q[4][0] ), .B(data_in[0]), .S(\wren[4] ), .Z(
        \din[4][0] ) );
    MUX21H MX1_1_4 ( .A(\q[4][1] ), .B(data_in[1]), .S(\wren[4] ), .Z(
        \din[4][1] ) );
    MUX21H MX1_1_14 ( .A(\q[14][1] ), .B(data_in[1]), .S(\wren[14] ), .Z(
        \din[14][1] ) );
    MUX21H MX1_2_8 ( .A(\q[8][2] ), .B(data_in[2]), .S(\wren[8] ), .Z(
        \din[8][2] ) );
    MUX21H MX1_0_5 ( .A(\q[5][0] ), .B(data_in[0]), .S(\wren[5] ), .Z(
        \din[5][0] ) );
    MUX21H MX1_0_14 ( .A(\q[14][0] ), .B(data_in[0]), .S(\wren[14] ), .Z(
        \din[14][0] ) );
    MUX21H MX1_0_15 ( .A(\q[15][0] ), .B(data_in[0]), .S(\wren[15] ), .Z(
        \din[15][0] ) );
    MUX21H MX1_5_2 ( .A(\q[2][5] ), .B(data_in[5]), .S(\wren[2] ), .Z(
        \din[2][5] ) );
    MUX21H MX1_6_10 ( .A(\q[10][6] ), .B(data_in[6]), .S(\wren[10] ), .Z(
        \din[10][6] ) );
    MUX21H MX1_8_5 ( .A(\q[5][8] ), .B(data_in[8]), .S(\wren[5] ), .Z(
        \din[5][8] ) );
    MUX21H MX1_12_7 ( .A(\q[7][12] ), .B(data_in[12]), .S(\wren[7] ), .Z(
        \din[7][12] ) );
    MUX21H MX1_12_13 ( .A(\q[13][12] ), .B(data_in[12]), .S(\wren[13] ), .Z(
        \din[13][12] ) );
    MUX21H MX1_2_0 ( .A(\q[0][2] ), .B(data_in[2]), .S(\wren[0] ), .Z(
        \din[0][2] ) );
    MUX21H MX1_2_10 ( .A(\q[10][2] ), .B(data_in[2]), .S(\wren[10] ), .Z(
        \din[10][2] ) );
    MUX21H MX1_4_15 ( .A(\q[15][4] ), .B(data_in[4]), .S(\wren[15] ), .Z(
        \din[15][4] ) );
    MUX21H MX1_10_3 ( .A(\q[3][10] ), .B(data_in[10]), .S(\wren[3] ), .Z(
        \din[3][10] ) );
    MUX21H MX1_15_5 ( .A(\q[5][15] ), .B(data_in[15]), .S(\wren[5] ), .Z(
        \din[5][15] ) );
    MUX21H MX1_3_0 ( .A(\q[0][3] ), .B(data_in[3]), .S(\wren[0] ), .Z(
        \din[0][3] ) );
    MUX21H MX1_5_14 ( .A(\q[14][5] ), .B(data_in[5]), .S(\wren[14] ), .Z(
        \din[14][5] ) );
    MUX21H MX1_6_6 ( .A(\q[6][6] ), .B(data_in[6]), .S(\wren[6] ), .Z(
        \din[6][6] ) );
    MUX21H MX1_7_6 ( .A(\q[6][7] ), .B(data_in[7]), .S(\wren[6] ), .Z(
        \din[6][7] ) );
    MUX21H MX1_3_11 ( .A(\q[11][3] ), .B(data_in[3]), .S(\wren[11] ), .Z(
        \din[11][3] ) );
    MUX21H MX1_11_3 ( .A(\q[3][11] ), .B(data_in[11]), .S(\wren[3] ), .Z(
        \din[3][11] ) );
    MUX21H MX1_12_6 ( .A(\q[6][12] ), .B(data_in[12]), .S(\wren[6] ), .Z(
        \din[6][12] ) );
    MUX21H MX1_14_5 ( .A(\q[5][14] ), .B(data_in[14]), .S(\wren[5] ), .Z(
        \din[5][14] ) );
    MUX21H MX1_8_4 ( .A(\q[4][8] ), .B(data_in[8]), .S(\wren[4] ), .Z(
        \din[4][8] ) );
    MUX21H MX1_12_12 ( .A(\q[12][12] ), .B(data_in[12]), .S(\wren[12] ), .Z(
        \din[12][12] ) );
    MUX21H MX1_2_9 ( .A(\q[9][2] ), .B(data_in[2]), .S(\wren[9] ), .Z(
        \din[9][2] ) );
    MUX21H MX1_3_9 ( .A(\q[9][3] ), .B(data_in[3]), .S(\wren[9] ), .Z(
        \din[9][3] ) );
    MUX21H MX1_5_3 ( .A(\q[3][5] ), .B(data_in[5]), .S(\wren[3] ), .Z(
        \din[3][5] ) );
    MUX21H MX1_6_11 ( .A(\q[11][6] ), .B(data_in[6]), .S(\wren[11] ), .Z(
        \din[11][6] ) );
    MUX21H MX1_4_3 ( .A(\q[3][4] ), .B(data_in[4]), .S(\wren[3] ), .Z(
        \din[3][4] ) );
    MUX21H MX1_13_13 ( .A(\q[13][13] ), .B(data_in[13]), .S(\wren[13] ), .Z(
        \din[13][13] ) );
    MUX21H MX1_1_2 ( .A(\q[2][1] ), .B(data_in[1]), .S(\wren[2] ), .Z(
        \din[2][1] ) );
    MUX21H MX1_1_5 ( .A(\q[5][1] ), .B(data_in[1]), .S(\wren[5] ), .Z(
        \din[5][1] ) );
    MUX21H MX1_1_12 ( .A(\q[12][1] ), .B(data_in[1]), .S(\wren[12] ), .Z(
        \din[12][1] ) );
    MUX21H MX1_1_15 ( .A(\q[15][1] ), .B(data_in[1]), .S(\wren[15] ), .Z(
        \din[15][1] ) );
    MUX21H MX1_6_8 ( .A(\q[8][6] ), .B(data_in[6]), .S(\wren[8] ), .Z(
        \din[8][6] ) );
    MUX21H MX1_13_6 ( .A(\q[6][13] ), .B(data_in[13]), .S(\wren[6] ), .Z(
        \din[6][13] ) );
    MUX21H MX1_7_10 ( .A(\q[10][7] ), .B(data_in[7]), .S(\wren[10] ), .Z(
        \din[10][7] ) );
    MUX21H MX1_9_3 ( .A(\q[3][9] ), .B(data_in[9]), .S(\wren[3] ), .Z(
        \din[3][9] ) );
    MUX21H MX1_9_4 ( .A(\q[4][9] ), .B(data_in[9]), .S(\wren[4] ), .Z(
        \din[4][9] ) );
    MUX21H MX1_13_1 ( .A(\q[1][13] ), .B(data_in[13]), .S(\wren[1] ), .Z(
        \din[1][13] ) );
    MUX21H MX1_15_11 ( .A(\q[11][15] ), .B(data_in[15]), .S(\wren[11] ), .Z(
        \din[11][15] ) );
    MUX21H MX1_4_4 ( .A(\q[4][4] ), .B(data_in[4]), .S(\wren[4] ), .Z(
        \din[4][4] ) );
    MUX21H MX1_13_14 ( .A(\q[14][13] ), .B(data_in[13]), .S(\wren[14] ), .Z(
        \din[14][13] ) );
    MUX21H MX1_7_8 ( .A(\q[8][7] ), .B(data_in[7]), .S(\wren[8] ), .Z(
        \din[8][7] ) );
    MUX21H MX1_5_4 ( .A(\q[4][5] ), .B(data_in[5]), .S(\wren[4] ), .Z(
        \din[4][5] ) );
    MUX21H MX1_14_10 ( .A(\q[10][14] ), .B(data_in[14]), .S(\wren[10] ), .Z(
        \din[10][14] ) );
    MUX21H MX1_0_13 ( .A(\q[13][0] ), .B(data_in[0]), .S(\wren[13] ), .Z(
        \din[13][0] ) );
    MUX21H MX1_12_1 ( .A(\q[1][12] ), .B(data_in[12]), .S(\wren[1] ), .Z(
        \din[1][12] ) );
    MUX21H MX1_8_3 ( .A(\q[3][8] ), .B(data_in[8]), .S(\wren[3] ), .Z(
        \din[3][8] ) );
    MUX21H MX1_9_10 ( .A(\q[10][9] ), .B(data_in[9]), .S(\wren[10] ), .Z(
        \din[10][9] ) );
    MUX21H MX1_11_10 ( .A(\q[10][11] ), .B(data_in[11]), .S(\wren[10] ), .Z(
        \din[10][11] ) );
    MUX21H MX1_12_15 ( .A(\q[15][12] ), .B(data_in[12]), .S(\wren[15] ), .Z(
        \din[15][12] ) );
    MUX21H MX1_13_8 ( .A(\q[8][13] ), .B(data_in[13]), .S(\wren[8] ), .Z(
        \din[8][13] ) );
    MUX21H MX1_14_2 ( .A(\q[2][14] ), .B(data_in[14]), .S(\wren[2] ), .Z(
        \din[2][14] ) );
    MUX21H MX1_11_4 ( .A(\q[4][11] ), .B(data_in[11]), .S(\wren[4] ), .Z(
        \din[4][11] ) );
    MUX21H MX1_2_7 ( .A(\q[7][2] ), .B(data_in[2]), .S(\wren[7] ), .Z(
        \din[7][2] ) );
    MUX21H MX1_3_7 ( .A(\q[7][3] ), .B(data_in[3]), .S(\wren[7] ), .Z(
        \din[7][3] ) );
    MUX21H MX1_5_13 ( .A(\q[13][5] ), .B(data_in[5]), .S(\wren[13] ), .Z(
        \din[13][5] ) );
    MUX21H MX1_6_1 ( .A(\q[1][6] ), .B(data_in[6]), .S(\wren[1] ), .Z(
        \din[1][6] ) );
    MUX21H MX1_7_1 ( .A(\q[1][7] ), .B(data_in[7]), .S(\wren[1] ), .Z(
        \din[1][7] ) );
    MUX21H MX1_10_11 ( .A(\q[11][10] ), .B(data_in[10]), .S(\wren[11] ), .Z(
        \din[11][10] ) );
    MUX21H MX1_4_12 ( .A(\q[12][4] ), .B(data_in[4]), .S(\wren[12] ), .Z(
        \din[12][4] ) );
    MUX21H MX1_8_11 ( .A(\q[11][8] ), .B(data_in[8]), .S(\wren[11] ), .Z(
        \din[11][8] ) );
    MUX21H MX1_12_8 ( .A(\q[8][12] ), .B(data_in[12]), .S(\wren[8] ), .Z(
        \din[8][12] ) );
    MUX21H MX1_10_4 ( .A(\q[4][10] ), .B(data_in[10]), .S(\wren[4] ), .Z(
        \din[4][10] ) );
    MUX21H MX1_15_2 ( .A(\q[2][15] ), .B(data_in[15]), .S(\wren[2] ), .Z(
        \din[2][15] ) );
    LD1 F0_11_13 ( .D(\din[13][11] ), .G(n38), .Q(\q[13][11] ) );
    LD1 F0_14_2 ( .D(\din[2][14] ), .G(n38), .Q(\q[2][14] ) );
    LD1 F0_9_10 ( .D(\din[10][9] ), .G(n38), .Q(\q[10][9] ) );
    LD1 F0_11_4 ( .D(\din[4][11] ), .G(n38), .Q(\q[4][11] ) );
    LD1 F0_5_13 ( .D(\din[13][5] ), .G(n38), .Q(\q[13][5] ) );
    LD1 F0_3_0 ( .D(\din[0][3] ), .G(n38), .Q(\q[0][3] ) );
    LD1 F0_13_8 ( .D(\din[8][13] ), .G(n38), .Q(\q[8][13] ) );
    LD1 F0_15_2 ( .D(\din[2][15] ), .G(n38), .Q(\q[2][15] ) );
    LD1 F0_10_4 ( .D(\din[4][10] ), .G(n38), .Q(\q[4][10] ) );
    LD1 F0_6_6 ( .D(\din[6][6] ), .G(n38), .Q(\q[6][6] ) );
    LD1 F0_10_12 ( .D(\din[12][10] ), .G(n38), .Q(\q[12][10] ) );
    LD1 F0_7_6 ( .D(\din[6][7] ), .G(n38), .Q(\q[6][7] ) );
    LD1 F0_12_8 ( .D(\din[8][12] ), .G(n38), .Q(\q[8][12] ) );
    LD1 F0_8_11 ( .D(\din[11][8] ), .G(n38), .Q(\q[11][8] ) );
    LD1 F0_4_12 ( .D(\din[12][4] ), .G(n38), .Q(\q[12][4] ) );
    LD1 F0_2_0 ( .D(\din[0][2] ), .G(n38), .Q(\q[0][2] ) );
    LD1 F0_9_4 ( .D(\din[4][9] ), .G(n38), .Q(\q[4][9] ) );
    LD1 F0_1_12 ( .D(\din[12][1] ), .G(n38), .Q(\q[12][1] ) );
    LD1 F0_15_12 ( .D(\din[12][15] ), .G(n38), .Q(\q[12][15] ) );
    LD1 F0_13_1 ( .D(\din[1][13] ), .G(n38), .Q(\q[1][13] ) );
    LD1 F0_4_3 ( .D(\din[3][4] ), .G(n38), .Q(\q[3][4] ) );
    LD1 F0_5_3 ( .D(\din[3][5] ), .G(n38), .Q(\q[3][5] ) );
    LD1 F0_3_9 ( .D(\din[9][3] ), .G(n38), .Q(\q[9][3] ) );
    LD1 F0_1_5 ( .D(\din[5][1] ), .G(n38), .Q(\q[5][1] ) );
    LD1 F0_0_13 ( .D(\din[13][0] ), .G(n38), .Q(\q[13][0] ) );
    LD1 F0_14_13 ( .D(\din[13][14] ), .G(n38), .Q(\q[13][14] ) );
    LD1 F0_12_1 ( .D(\din[1][12] ), .G(n38), .Q(\q[1][12] ) );
    LD1 F0_8_4 ( .D(\din[4][8] ), .G(n38), .Q(\q[4][8] ) );
    LD1 F0_12_11 ( .D(\din[11][12] ), .G(n38), .Q(\q[11][12] ) );
    LD1 F0_8_3 ( .D(\din[3][8] ), .G(n38), .Q(\q[3][8] ) );
    LD1 F0_6_11 ( .D(\din[11][6] ), .G(n38), .Q(\q[11][6] ) );
    LD1 F0_2_9 ( .D(\din[9][2] ), .G(n38), .Q(\q[9][2] ) );
    LD1 F0_14_14 ( .D(\din[14][14] ), .G(n38), .Q(\q[14][14] ) );
    LD1 F0_0_5 ( .D(\din[5][0] ), .G(n38), .Q(\q[5][0] ) );
    LD1 F0_7_8 ( .D(\din[8][7] ), .G(n38), .Q(\q[8][7] ) );
    LD1 F0_5_4 ( .D(\din[4][5] ), .G(n38), .Q(\q[4][5] ) );
    LD1 F0_13_10 ( .D(\din[10][13] ), .G(n38), .Q(\q[10][13] ) );
    LD1 F0_12_6 ( .D(\din[6][12] ), .G(n38), .Q(\q[6][12] ) );
    LD1 F0_4_4 ( .D(\din[4][4] ), .G(n38), .Q(\q[4][4] ) );
    LD1 F0_7_10 ( .D(\din[10][7] ), .G(n38), .Q(\q[10][7] ) );
    LD1 F0_1_2 ( .D(\din[2][1] ), .G(n38), .Q(\q[2][1] ) );
    LD1 F0_0_14 ( .D(\din[14][0] ), .G(n38), .Q(\q[14][0] ) );
    LD1 F0_13_6 ( .D(\din[6][13] ), .G(n38), .Q(\q[6][13] ) );
    LD1 F0_15_15 ( .D(\din[15][15] ), .G(n38), .Q(\q[15][15] ) );
    LD1 F0_6_8 ( .D(\din[8][6] ), .G(n38), .Q(\q[8][6] ) );
    LD1 F0_9_3 ( .D(\din[3][9] ), .G(n38), .Q(\q[3][9] ) );
    LD1 F0_15_5 ( .D(\din[5][15] ), .G(n38), .Q(\q[5][15] ) );
    LD1 F0_10_3 ( .D(\din[3][10] ), .G(n38), .Q(\q[3][10] ) );
    LD1 F0_4_15 ( .D(\din[15][4] ), .G(n38), .Q(\q[15][4] ) );
    LD1 F0_2_10 ( .D(\din[10][2] ), .G(n38), .Q(\q[10][2] ) );
    LD1 F0_10_15 ( .D(\din[15][10] ), .G(n38), .Q(\q[15][10] ) );
    LD1 F0_7_1 ( .D(\din[1][7] ), .G(n38), .Q(\q[1][7] ) );
    LD1 F0_14_5 ( .D(\din[5][14] ), .G(n38), .Q(\q[5][14] ) );
    LD1 F0_11_3 ( .D(\din[3][11] ), .G(n38), .Q(\q[3][11] ) );
    LD1 F0_6_1 ( .D(\din[1][6] ), .G(n38), .Q(\q[1][6] ) );
    LD1 F0_3_11 ( .D(\din[11][3] ), .G(n38), .Q(\q[11][3] ) );
    LD1 F0_2_7 ( .D(\din[7][2] ), .G(n38), .Q(\q[7][2] ) );
    LD1 F0_11_14 ( .D(\din[14][11] ), .G(n38), .Q(\q[14][11] ) );
    LD1 F0_5_14 ( .D(\din[14][5] ), .G(n38), .Q(\q[14][5] ) );
    LD1 F0_15_14 ( .D(\din[14][15] ), .G(n38), .Q(\q[14][15] ) );
    LD1 F0_3_7 ( .D(\din[7][3] ), .G(n38), .Q(\q[7][3] ) );
    LD1 F0_1_15 ( .D(\din[15][1] ), .G(n38), .Q(\q[15][1] ) );
    LD1 F0_9_2 ( .D(\din[2][9] ), .G(n38), .Q(\q[2][9] ) );
    LD1 F0_13_11 ( .D(\din[11][13] ), .G(n38), .Q(\q[11][13] ) );
    LD1 F0_4_5 ( .D(\din[5][4] ), .G(n38), .Q(\q[5][4] ) );
    LD1 F0_1_14 ( .D(\din[14][1] ), .G(n38), .Q(\q[14][1] ) );
    LD1 F0_1_3 ( .D(\din[3][1] ), .G(n38), .Q(\q[3][1] ) );
    LD1 F0_13_7 ( .D(\din[7][13] ), .G(n38), .Q(\q[7][13] ) );
    LD1 F0_7_11 ( .D(\din[11][7] ), .G(n38), .Q(\q[11][7] ) );
    LD1 F0_6_9 ( .D(\din[9][6] ), .G(n38), .Q(\q[9][6] ) );
    LD1 F0_14_15 ( .D(\din[15][14] ), .G(n38), .Q(\q[15][14] ) );
    LD1 F0_12_7 ( .D(\din[7][12] ), .G(n38), .Q(\q[7][12] ) );
    LD1 F0_7_9 ( .D(\din[9][7] ), .G(n38), .Q(\q[9][7] ) );
    LD1 F0_5_5 ( .D(\din[5][5] ), .G(n38), .Q(\q[5][5] ) );
    LD1 F0_12_10 ( .D(\din[10][12] ), .G(n38), .Q(\q[10][12] ) );
    LD1 F0_8_2 ( .D(\din[2][8] ), .G(n38), .Q(\q[2][8] ) );
    LD1 F0_6_10 ( .D(\din[10][6] ), .G(n38), .Q(\q[10][6] ) );
    LD1 F0_11_15 ( .D(\din[15][11] ), .G(n38), .Q(\q[15][11] ) );
    LD1 F0_5_15 ( .D(\din[15][5] ), .G(n38), .Q(\q[15][5] ) );
    LD1 F0_14_4 ( .D(\din[4][14] ), .G(n38), .Q(\q[4][14] ) );
    LD1 F0_11_2 ( .D(\din[2][11] ), .G(n38), .Q(\q[2][11] ) );
    LD1 F0_6_0 ( .D(\din[0][6] ), .G(n38), .Q(\q[0][6] ) );
    LD1 F0_3_10 ( .D(\din[10][3] ), .G(n38), .Q(\q[10][3] ) );
    LD1 F0_3_6 ( .D(\din[6][3] ), .G(n38), .Q(\q[6][3] ) );
    LD1 F0_15_4 ( .D(\din[4][15] ), .G(n38), .Q(\q[4][15] ) );
    LD1 F0_10_2 ( .D(\din[2][10] ), .G(n38), .Q(\q[2][10] ) );
    LD1 F0_4_14 ( .D(\din[14][4] ), .G(n38), .Q(\q[14][4] ) );
    LD1 F0_7_0 ( .D(\din[0][7] ), .G(n38), .Q(\q[0][7] ) );
    LD1 F0_10_14 ( .D(\din[14][10] ), .G(n38), .Q(\q[14][10] ) );
    LD1 F0_15_3 ( .D(\din[3][15] ), .G(n38), .Q(\q[3][15] ) );
    LD1 F0_10_13 ( .D(\din[13][10] ), .G(n38), .Q(\q[13][10] ) );
    LD1 F0_10_5 ( .D(\din[5][10] ), .G(n38), .Q(\q[5][10] ) );
    LD1 F0_8_10 ( .D(\din[10][8] ), .G(n38), .Q(\q[10][8] ) );
    LD1 F0_12_9 ( .D(\din[9][12] ), .G(n38), .Q(\q[9][12] ) );
    LD1 F0_7_7 ( .D(\din[7][7] ), .G(n38), .Q(\q[7][7] ) );
    LD1 F0_2_11 ( .D(\din[11][2] ), .G(n38), .Q(\q[11][2] ) );
    LD1 F0_2_6 ( .D(\din[6][2] ), .G(n38), .Q(\q[6][2] ) );
    LD1 F0_14_3 ( .D(\din[3][14] ), .G(n38), .Q(\q[3][14] ) );
    LD1 F0_9_11 ( .D(\din[11][9] ), .G(n38), .Q(\q[11][9] ) );
    LD1 F0_11_5 ( .D(\din[5][11] ), .G(n38), .Q(\q[5][11] ) );
    LD1 F0_4_13 ( .D(\din[13][4] ), .G(n38), .Q(\q[13][4] ) );
    LD1 F0_13_9 ( .D(\din[9][13] ), .G(n38), .Q(\q[9][13] ) );
    LD1 F0_3_1 ( .D(\din[1][3] ), .G(n38), .Q(\q[1][3] ) );
    LD1 F0_6_7 ( .D(\din[7][6] ), .G(n38), .Q(\q[7][6] ) );
    LD1 F0_11_12 ( .D(\din[12][11] ), .G(n38), .Q(\q[12][11] ) );
    LD1 F0_8_5 ( .D(\din[5][8] ), .G(n38), .Q(\q[5][8] ) );
    LD1 F0_5_12 ( .D(\din[12][5] ), .G(n38), .Q(\q[12][5] ) );
    LD1 F0_5_2 ( .D(\din[2][5] ), .G(n38), .Q(\q[2][5] ) );
    LD1 F0_2_1 ( .D(\din[1][2] ), .G(n38), .Q(\q[1][2] ) );
    LD1 F0_0_15 ( .D(\din[15][0] ), .G(n38), .Q(\q[15][0] ) );
    LD1 F0_14_12 ( .D(\din[12][14] ), .G(n38), .Q(\q[12][14] ) );
    LD1 F0_0_12 ( .D(\din[12][0] ), .G(n38), .Q(\q[12][0] ) );
    LD1 F0_12_0 ( .D(\din[0][12] ), .G(n38), .Q(\q[0][12] ) );
    LD1 F0_2_8 ( .D(\din[8][2] ), .G(n38), .Q(\q[8][2] ) );
    LD1 F0_0_4 ( .D(\din[4][0] ), .G(n38), .Q(\q[4][0] ) );
    LD1 F0_0_3 ( .D(\din[3][0] ), .G(n38), .Q(\q[3][0] ) );
    LD1 F0_13_0 ( .D(\din[0][13] ), .G(n38), .Q(\q[0][13] ) );
    LD1 F0_4_2 ( .D(\din[2][4] ), .G(n38), .Q(\q[2][4] ) );
    LD1 F0_3_8 ( .D(\din[8][3] ), .G(n38), .Q(\q[8][3] ) );
    LD1 F0_9_5 ( .D(\din[5][9] ), .G(n38), .Q(\q[5][9] ) );
    LD1 F0_1_13 ( .D(\din[13][1] ), .G(n38), .Q(\q[13][1] ) );
    LD1 F0_1_4 ( .D(\din[4][1] ), .G(n38), .Q(\q[4][1] ) );
    LD1 F0_15_13 ( .D(\din[13][15] ), .G(n38), .Q(\q[13][15] ) );
    LD1 F0_5_10 ( .D(\din[10][5] ), .G(n38), .Q(\q[10][5] ) );
    LD1 F0_11_10 ( .D(\din[10][11] ), .G(n38), .Q(\q[10][11] ) );
    LD1 F0_6_5 ( .D(\din[5][6] ), .G(n38), .Q(\q[5][6] ) );
    LD1 F0_3_15 ( .D(\din[15][3] ), .G(n38), .Q(\q[15][3] ) );
    LD1 F0_3_3 ( .D(\din[3][3] ), .G(n38), .Q(\q[3][3] ) );
    LD1 F0_11_7 ( .D(\din[7][11] ), .G(n38), .Q(\q[7][11] ) );
    LD1 F0_9_13 ( .D(\din[13][9] ), .G(n38), .Q(\q[13][9] ) );
    LD1 F0_14_1 ( .D(\din[1][14] ), .G(n38), .Q(\q[1][14] ) );
    LD1 F0_4_9 ( .D(\din[9][4] ), .G(n38), .Q(\q[9][4] ) );
    LD1 F0_4_11 ( .D(\din[11][4] ), .G(n38), .Q(\q[11][4] ) );
    LD1 F0_10_11 ( .D(\din[11][10] ), .G(n38), .Q(\q[11][10] ) );
    LD1 F0_7_5 ( .D(\din[5][7] ), .G(n38), .Q(\q[5][7] ) );
    LD1 F0_15_1 ( .D(\din[1][15] ), .G(n38), .Q(\q[1][15] ) );
    LD1 F0_10_7 ( .D(\din[7][10] ), .G(n38), .Q(\q[7][10] ) );
    LD1 F0_5_9 ( .D(\din[9][5] ), .G(n38), .Q(\q[9][5] ) );
    LD1 F0_2_3 ( .D(\din[3][2] ), .G(n38), .Q(\q[3][2] ) );
    LD1 F0_8_12 ( .D(\din[12][8] ), .G(n38), .Q(\q[12][8] ) );
    LD1 F0_2_14 ( .D(\din[14][2] ), .G(n38), .Q(\q[14][2] ) );
    LD1 F0_15_11 ( .D(\din[11][15] ), .G(n38), .Q(\q[11][15] ) );
    LD1 F0_13_2 ( .D(\din[2][13] ), .G(n38), .Q(\q[2][13] ) );
    LD1 F0_9_7 ( .D(\din[7][9] ), .G(n38), .Q(\q[7][9] ) );
    LD1 F0_14_8 ( .D(\din[8][14] ), .G(n38), .Q(\q[8][14] ) );
    LD1 F0_13_14 ( .D(\din[14][13] ), .G(n38), .Q(\q[14][13] ) );
    LD1 F0_4_0 ( .D(\din[0][4] ), .G(n38), .Q(\q[0][4] ) );
    LD1 F0_1_11 ( .D(\din[11][1] ), .G(n38), .Q(\q[11][1] ) );
    LD1 F0_0_2 ( .D(\din[2][0] ), .G(n38), .Q(\q[2][0] ) );
    LD1 F0_7_14 ( .D(\din[14][7] ), .G(n38), .Q(\q[14][7] ) );
    LD1 F0_12_2 ( .D(\din[2][12] ), .G(n38), .Q(\q[2][12] ) );
    LD1 F0_1_6 ( .D(\din[6][1] ), .G(n38), .Q(\q[6][1] ) );
    LD1 F0_14_10 ( .D(\din[10][14] ), .G(n38), .Q(\q[10][14] ) );
    LD1 F0_5_0 ( .D(\din[0][5] ), .G(n38), .Q(\q[0][5] ) );
    LD1 F0_15_8 ( .D(\din[8][15] ), .G(n38), .Q(\q[8][15] ) );
    LD1 F0_12_15 ( .D(\din[15][12] ), .G(n38), .Q(\q[15][12] ) );
    LD1 F0_8_7 ( .D(\din[7][8] ), .G(n38), .Q(\q[7][8] ) );
    LD1 F0_6_15 ( .D(\din[15][6] ), .G(n38), .Q(\q[15][6] ) );
    LD1 F0_12_12 ( .D(\din[12][12] ), .G(n38), .Q(\q[12][12] ) );
    LD1 F0_12_5 ( .D(\din[5][12] ), .G(n38), .Q(\q[5][12] ) );
    LD1 F0_8_0 ( .D(\din[0][8] ), .G(n38), .Q(\q[0][8] ) );
    LD1 F0_6_12 ( .D(\din[12][6] ), .G(n38), .Q(\q[12][6] ) );
    LD1 F0_10_9 ( .D(\din[9][10] ), .G(n38), .Q(\q[9][10] ) );
    LD1 F0_5_7 ( .D(\din[7][5] ), .G(n38), .Q(\q[7][5] ) );
    LD1 F0_0_10 ( .D(\din[10][0] ), .G(n38), .Q(\q[10][0] ) );
    LD1 F0_0_6 ( .D(\din[6][0] ), .G(n38), .Q(\q[6][0] ) );
    LD1 F0_13_5 ( .D(\din[5][13] ), .G(n38), .Q(\q[5][13] ) );
    LD1 F0_11_9 ( .D(\din[9][11] ), .G(n38), .Q(\q[9][11] ) );
    LD1 F0_7_13 ( .D(\din[13][7] ), .G(n38), .Q(\q[13][7] ) );
    LD1 F0_1_1 ( .D(\din[1][1] ), .G(n38), .Q(\q[1][1] ) );
    LD1 F0_13_13 ( .D(\din[13][13] ), .G(n38), .Q(\q[13][13] ) );
    LD1 F0_9_0 ( .D(\din[0][9] ), .G(n38), .Q(\q[0][9] ) );
    LD1 F0_4_7 ( .D(\din[7][4] ), .G(n38), .Q(\q[7][4] ) );
    LD1 F0_8_15 ( .D(\din[15][8] ), .G(n38), .Q(\q[15][8] ) );
    LD1 F0_8_9 ( .D(\din[9][8] ), .G(n38), .Q(\q[9][8] ) );
    LD1 F0_7_2 ( .D(\din[2][7] ), .G(n38), .Q(\q[2][7] ) );
    LD1 F0_2_13 ( .D(\din[13][2] ), .G(n38), .Q(\q[13][2] ) );
    LD1 F0_2_4 ( .D(\din[4][2] ), .G(n38), .Q(\q[4][2] ) );
    LD1 F0_10_0 ( .D(\din[0][10] ), .G(n38), .Q(\q[0][10] ) );
    LD1 F0_15_6 ( .D(\din[6][15] ), .G(n38), .Q(\q[6][15] ) );
    LD1 F0_3_4 ( .D(\din[4][3] ), .G(n38), .Q(\q[4][3] ) );
    LD1 F0_6_2 ( .D(\din[2][6] ), .G(n38), .Q(\q[2][6] ) );
    LD1 F0_14_6 ( .D(\din[6][14] ), .G(n38), .Q(\q[6][14] ) );
    LD1 F0_11_0 ( .D(\din[0][11] ), .G(n38), .Q(\q[0][11] ) );
    LD1 F0_9_14 ( .D(\din[14][9] ), .G(n38), .Q(\q[14][9] ) );
    LD1 F0_3_12 ( .D(\din[12][3] ), .G(n38), .Q(\q[12][3] ) );
    LD1 F0_9_9 ( .D(\din[9][9] ), .G(n38), .Q(\q[9][9] ) );
    LD1 F0_9_1 ( .D(\din[1][9] ), .G(n38), .Q(\q[1][9] ) );
    LD1 F0_13_4 ( .D(\din[4][13] ), .G(n38), .Q(\q[4][13] ) );
    LD1 F0_1_8 ( .D(\din[8][1] ), .G(n38), .Q(\q[8][1] ) );
    LD1 F0_1_0 ( .D(\din[0][1] ), .G(n38), .Q(\q[0][1] ) );
    LD1 F0_0_8 ( .D(\din[8][0] ), .G(n38), .Q(\q[8][0] ) );
    LD1 F0_11_8 ( .D(\din[8][11] ), .G(n38), .Q(\q[8][11] ) );
    LD1 F0_13_12 ( .D(\din[12][13] ), .G(n38), .Q(\q[12][13] ) );
    LD1 F0_7_12 ( .D(\din[12][7] ), .G(n38), .Q(\q[12][7] ) );
    LD1 F0_12_4 ( .D(\din[4][12] ), .G(n38), .Q(\q[4][12] ) );
    LD1 F0_4_6 ( .D(\din[6][4] ), .G(n38), .Q(\q[6][4] ) );
    LD1 F0_5_6 ( .D(\din[6][5] ), .G(n38), .Q(\q[6][5] ) );
    LD1 F0_10_8 ( .D(\din[8][10] ), .G(n38), .Q(\q[8][10] ) );
    LD1 F0_0_1 ( .D(\din[1][0] ), .G(n38), .Q(\q[1][0] ) );
    LD1 F0_12_13 ( .D(\din[13][12] ), .G(n38), .Q(\q[13][12] ) );
    LD1 F0_9_8 ( .D(\din[8][9] ), .G(n38), .Q(\q[8][9] ) );
    LD1 F0_8_1 ( .D(\din[1][8] ), .G(n38), .Q(\q[1][8] ) );
    LD1 F0_6_13 ( .D(\din[13][6] ), .G(n38), .Q(\q[13][6] ) );
    LD1 F0_6_3 ( .D(\din[3][6] ), .G(n38), .Q(\q[3][6] ) );
    LD1 F0_14_7 ( .D(\din[7][14] ), .G(n38), .Q(\q[7][14] ) );
    LD1 F0_11_1 ( .D(\din[1][11] ), .G(n38), .Q(\q[1][11] ) );
    LD1 F0_9_15 ( .D(\din[15][9] ), .G(n38), .Q(\q[15][9] ) );
    LD1 F0_3_13 ( .D(\din[13][3] ), .G(n38), .Q(\q[13][3] ) );
    LD1 F0_3_5 ( .D(\din[5][3] ), .G(n38), .Q(\q[5][3] ) );
    LD1 F0_7_3 ( .D(\din[3][7] ), .G(n38), .Q(\q[3][7] ) );
    LD1 F0_2_5 ( .D(\din[5][2] ), .G(n38), .Q(\q[5][2] ) );
    LD1 F0_1_9 ( .D(\din[9][1] ), .G(n38), .Q(\q[9][1] ) );
    LD1 F0_15_7 ( .D(\din[7][15] ), .G(n38), .Q(\q[7][15] ) );
    LD1 F0_10_1 ( .D(\din[1][10] ), .G(n38), .Q(\q[1][10] ) );
    LD1 F0_8_14 ( .D(\din[14][8] ), .G(n38), .Q(\q[14][8] ) );
    LD1 F0_8_8 ( .D(\din[8][8] ), .G(n38), .Q(\q[8][8] ) );
    LD1 F0_8_13 ( .D(\din[13][8] ), .G(n38), .Q(\q[13][8] ) );
    LD1 F0_4_10 ( .D(\din[10][4] ), .G(n38), .Q(\q[10][4] ) );
    LD1 F0_2_15 ( .D(\din[15][2] ), .G(n38), .Q(\q[15][2] ) );
    LD1 F0_2_12 ( .D(\din[12][2] ), .G(n38), .Q(\q[12][2] ) );
    LD1 F0_10_10 ( .D(\din[10][10] ), .G(n38), .Q(\q[10][10] ) );
    LD1 F0_15_0 ( .D(\din[0][15] ), .G(n38), .Q(\q[0][15] ) );
    LD1 F0_7_4 ( .D(\din[4][7] ), .G(n38), .Q(\q[4][7] ) );
    LD1 F0_5_8 ( .D(\din[8][5] ), .G(n38), .Q(\q[8][5] ) );
    LD1 F0_2_2 ( .D(\din[2][2] ), .G(n38), .Q(\q[2][2] ) );
    LD1 F0_10_6 ( .D(\din[6][10] ), .G(n38), .Q(\q[6][10] ) );
    LD1 F0_6_4 ( .D(\din[4][6] ), .G(n38), .Q(\q[4][6] ) );
    LD1 F0_3_14 ( .D(\din[14][3] ), .G(n38), .Q(\q[14][3] ) );
    LD1 F0_3_2 ( .D(\din[2][3] ), .G(n38), .Q(\q[2][3] ) );
    LD1 F0_0_9 ( .D(\din[9][0] ), .G(n38), .Q(\q[9][0] ) );
    LD1 F0_11_6 ( .D(\din[6][11] ), .G(n38), .Q(\q[6][11] ) );
    LD1 F0_14_0 ( .D(\din[0][14] ), .G(n38), .Q(\q[0][14] ) );
    LD1 F0_9_12 ( .D(\din[12][9] ), .G(n38), .Q(\q[12][9] ) );
    LD1 F0_5_11 ( .D(\din[11][5] ), .G(n38), .Q(\q[11][5] ) );
    LD1 F0_11_11 ( .D(\din[11][11] ), .G(n38), .Q(\q[11][11] ) );
    LD1 F0_12_14 ( .D(\din[14][12] ), .G(n38), .Q(\q[14][12] ) );
    LD1 F0_8_6 ( .D(\din[6][8] ), .G(n38), .Q(\q[6][8] ) );
    LD1 F0_14_11 ( .D(\din[11][14] ), .G(n38), .Q(\q[11][14] ) );
    LD1 F0_12_3 ( .D(\din[3][12] ), .G(n38), .Q(\q[3][12] ) );
    LD1 F0_6_14 ( .D(\din[14][6] ), .G(n38), .Q(\q[14][6] ) );
    LD1 F0_4_8 ( .D(\din[8][4] ), .G(n38), .Q(\q[8][4] ) );
    LD1 F0_15_9 ( .D(\din[9][15] ), .G(n38), .Q(\q[9][15] ) );
    LD1 F0_5_1 ( .D(\din[1][5] ), .G(n38), .Q(\q[1][5] ) );
    LD1 F0_14_9 ( .D(\din[9][14] ), .G(n38), .Q(\q[9][14] ) );
    LD1 F0_13_3 ( .D(\din[3][13] ), .G(n38), .Q(\q[3][13] ) );
    LD1 F0_13_15 ( .D(\din[15][13] ), .G(n38), .Q(\q[15][13] ) );
    LD1 F0_7_15 ( .D(\din[15][7] ), .G(n38), .Q(\q[15][7] ) );
    LD1 F0_4_1 ( .D(\din[1][4] ), .G(n38), .Q(\q[1][4] ) );
    LD1 F0_0_11 ( .D(\din[11][0] ), .G(n38), .Q(\q[11][0] ) );
    LD1 F0_0_7 ( .D(\din[7][0] ), .G(n38), .Q(\q[7][0] ) );
    LD1 F0_0_0 ( .D(\din[0][0] ), .G(n38), .Q(\q[0][0] ) );
    LD1 F0_1_7 ( .D(\din[7][1] ), .G(n38), .Q(\q[7][1] ) );
    LD1 F0_15_10 ( .D(\din[10][15] ), .G(n38), .Q(\q[10][15] ) );
    LD1 F0_9_6 ( .D(\din[6][9] ), .G(n38), .Q(\q[6][9] ) );
    LD1 F0_1_10 ( .D(\din[10][1] ), .G(n38), .Q(\q[10][1] ) );
    NR2 U39 ( .A(n39), .B(wr_n), .Z(\wren[6] ) );
    NR2 U40 ( .A(n40), .B(wr_n), .Z(\wren[1] ) );
    NR2 U41 ( .A(n41), .B(wr_n), .Z(\wren[8] ) );
    NR2 U42 ( .A(n42), .B(wr_n), .Z(\wren[10] ) );
    NR2 U43 ( .A(n43), .B(wr_n), .Z(\wren[0] ) );
    NR2 U44 ( .A(n44), .B(wr_n), .Z(\wren[11] ) );
    NR2 U45 ( .A(n45), .B(wr_n), .Z(\wren[9] ) );
    NR2 U46 ( .A(n46), .B(wr_n), .Z(\wren[7] ) );
    NR2 U47 ( .A(n47), .B(wr_n), .Z(\wren[14] ) );
    NR2 U48 ( .A(n48), .B(wr_n), .Z(\wren[5] ) );
    NR2 U49 ( .A(n49), .B(wr_n), .Z(\wren[2] ) );
    NR2 U50 ( .A(n50), .B(wr_n), .Z(\wren[13] ) );
    NR2 U51 ( .A(n51), .B(wr_n), .Z(\wren[3] ) );
    NR2 U52 ( .A(n52), .B(wr_n), .Z(\wren[12] ) );
    NR2 U53 ( .A(n53), .B(wr_n), .Z(\wren[15] ) );
    NR2 U54 ( .A(n54), .B(wr_n), .Z(\wren[4] ) );
    IV U55 ( .A(clk), .Z(n38) );
    IV U56 ( .A(wr_addr[9]), .Z(n45) );
    IV U57 ( .A(wr_addr[8]), .Z(n41) );
    IV U58 ( .A(wr_addr[7]), .Z(n46) );
    IV U59 ( .A(wr_addr[6]), .Z(n39) );
    IV U60 ( .A(wr_addr[5]), .Z(n48) );
    IV U61 ( .A(wr_addr[4]), .Z(n54) );
    IV U62 ( .A(wr_addr[3]), .Z(n51) );
    IV U63 ( .A(wr_addr[2]), .Z(n49) );
    IV U64 ( .A(wr_addr[1]), .Z(n40) );
    IV U65 ( .A(wr_addr[15]), .Z(n53) );
    IV U66 ( .A(wr_addr[14]), .Z(n47) );
    IV U67 ( .A(wr_addr[13]), .Z(n50) );
    IV U68 ( .A(wr_addr[12]), .Z(n52) );
    IV U69 ( .A(wr_addr[11]), .Z(n44) );
    IV U70 ( .A(wr_addr[10]), .Z(n42) );
    IV U71 ( .A(wr_addr[0]), .Z(n43) );
endmodule


module fifo_DW01_mux_any_256_4_16_0 ( A, SEL, MUX );
input  [255:0] A;
input  [3:0] SEL;
output [15:0] MUX;
    wire \tmp[3][136] , \tmp[3][14] , \tmp[3][132] , \tmp[3][10] , 
        \tmp[3][139] , \tmp[3][130] , \tmp[3][129] , \tmp[3][12] , 
        \tmp[3][134] , \tmp[3][1] , \tmp[3][8] , \tmp[3][141] , \tmp[3][5] , 
        \tmp[3][7] , \tmp[3][143] , \tmp[3][3] , \tmp[3][142] , \tmp[3][2] , 
        \tmp[3][6] , \tmp[3][4] , \tmp[3][0] , \tmp[3][9] , \tmp[3][140] , 
        \tmp[3][135] , \tmp[3][138] , \tmp[3][13] , \tmp[3][131] , 
        \tmp[3][128] , \tmp[3][11] , \tmp[3][133] , \tmp[3][137] , 
        \tmp[3][15] , n56, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, 
        n68, n69, n70, n71, n72, n73;
    MUX81P MX8_1_1_0 ( .D0(A[0]), .D1(A[16]), .D2(A[32]), .D3(A[48]), .D4(A
        [64]), .D5(A[80]), .D6(A[96]), .D7(A[112]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][0] ) );
    MUX81P MX8_1_1_1 ( .D0(A[1]), .D1(A[17]), .D2(A[33]), .D3(A[49]), .D4(A
        [65]), .D5(A[81]), .D6(A[97]), .D7(A[113]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][1] ) );
    MUX81P MX8_1_1_2 ( .D0(A[2]), .D1(A[18]), .D2(A[34]), .D3(A[50]), .D4(A
        [66]), .D5(A[82]), .D6(A[98]), .D7(A[114]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][2] ) );
    MUX81P MX8_1_5_10 ( .D0(A[138]), .D1(A[154]), .D2(A[170]), .D3(A[186]), 
        .D4(A[202]), .D5(A[218]), .D6(A[234]), .D7(A[250]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][138] ) );
    MUX81P MX8_1_1_3 ( .D0(A[3]), .D1(A[19]), .D2(A[35]), .D3(A[51]), .D4(A
        [67]), .D5(A[83]), .D6(A[99]), .D7(A[115]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][3] ) );
    MUX81P MX8_1_1_4 ( .D0(A[4]), .D1(A[20]), .D2(A[36]), .D3(A[52]), .D4(A
        [68]), .D5(A[84]), .D6(A[100]), .D7(A[116]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][4] ) );
    MUX81P MX8_1_1_5 ( .D0(A[5]), .D1(A[21]), .D2(A[37]), .D3(A[53]), .D4(A
        [69]), .D5(A[85]), .D6(A[101]), .D7(A[117]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][5] ) );
    MUX81P MX8_1_1_11 ( .D0(A[11]), .D1(A[27]), .D2(A[43]), .D3(A[59]), .D4(A
        [75]), .D5(A[91]), .D6(A[107]), .D7(A[123]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][11] ) );
    MUX81P MX8_1_5_3 ( .D0(A[131]), .D1(A[147]), .D2(A[163]), .D3(A[179]), 
        .D4(A[195]), .D5(A[211]), .D6(A[227]), .D7(A[243]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][131] ) );
    MUX81P MX8_1_5_4 ( .D0(A[132]), .D1(A[148]), .D2(A[164]), .D3(A[180]), 
        .D4(A[196]), .D5(A[212]), .D6(A[228]), .D7(A[244]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][132] ) );
    MUX81P MX8_1_1_10 ( .D0(A[10]), .D1(A[26]), .D2(A[42]), .D3(A[58]), .D4(A
        [74]), .D5(A[90]), .D6(A[106]), .D7(A[122]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][10] ) );
    MUX81P MX8_1_5_2 ( .D0(A[130]), .D1(A[146]), .D2(A[162]), .D3(A[178]), 
        .D4(A[194]), .D5(A[210]), .D6(A[226]), .D7(A[242]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][130] ) );
    MUX81P MX8_1_5_5 ( .D0(A[133]), .D1(A[149]), .D2(A[165]), .D3(A[181]), 
        .D4(A[197]), .D5(A[213]), .D6(A[229]), .D7(A[245]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][133] ) );
    MUX81P MX8_1_5_11 ( .D0(A[139]), .D1(A[155]), .D2(A[171]), .D3(A[187]), 
        .D4(A[203]), .D5(A[219]), .D6(A[235]), .D7(A[251]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][139] ) );
    MUX81P MX8_1_1_8 ( .D0(A[8]), .D1(A[24]), .D2(A[40]), .D3(A[56]), .D4(A
        [72]), .D5(A[88]), .D6(A[104]), .D7(A[120]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][8] ) );
    MUX81P MX8_1_5_13 ( .D0(A[141]), .D1(A[157]), .D2(A[173]), .D3(A[189]), 
        .D4(A[205]), .D5(A[221]), .D6(A[237]), .D7(A[253]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][141] ) );
    MUX81P MX8_1_1_6 ( .D0(A[6]), .D1(A[22]), .D2(A[38]), .D3(A[54]), .D4(A
        [70]), .D5(A[86]), .D6(A[102]), .D7(A[118]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][6] ) );
    MUX81P MX8_1_1_12 ( .D0(A[12]), .D1(A[28]), .D2(A[44]), .D3(A[60]), .D4(A
        [76]), .D5(A[92]), .D6(A[108]), .D7(A[124]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][12] ) );
    MUX81P MX8_1_1_15 ( .D0(A[15]), .D1(A[31]), .D2(A[47]), .D3(A[63]), .D4(A
        [79]), .D5(A[95]), .D6(A[111]), .D7(A[127]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][15] ) );
    MUX81P MX8_1_5_0 ( .D0(A[128]), .D1(A[144]), .D2(A[160]), .D3(A[176]), 
        .D4(A[192]), .D5(A[208]), .D6(A[224]), .D7(A[240]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][128] ) );
    MUX81P MX8_1_5_7 ( .D0(A[135]), .D1(A[151]), .D2(A[167]), .D3(A[183]), 
        .D4(A[199]), .D5(A[215]), .D6(A[231]), .D7(A[247]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][135] ) );
    MUX81P MX8_1_1_7 ( .D0(A[7]), .D1(A[23]), .D2(A[39]), .D3(A[55]), .D4(A
        [71]), .D5(A[87]), .D6(A[103]), .D7(A[119]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][7] ) );
    MUX81P MX8_1_5_9 ( .D0(A[137]), .D1(A[153]), .D2(A[169]), .D3(A[185]), 
        .D4(A[201]), .D5(A[217]), .D6(A[233]), .D7(A[249]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][137] ) );
    MUX81P MX8_1_5_14 ( .D0(A[142]), .D1(A[158]), .D2(A[174]), .D3(A[190]), 
        .D4(A[206]), .D5(A[222]), .D6(A[238]), .D7(A[254]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][142] ) );
    MUX81P MX8_1_1_9 ( .D0(A[9]), .D1(A[25]), .D2(A[41]), .D3(A[57]), .D4(A
        [73]), .D5(A[89]), .D6(A[105]), .D7(A[121]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][9] ) );
    MUX81P MX8_1_1_14 ( .D0(A[14]), .D1(A[30]), .D2(A[46]), .D3(A[62]), .D4(A
        [78]), .D5(A[94]), .D6(A[110]), .D7(A[126]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][14] ) );
    MUX81P MX8_1_5_1 ( .D0(A[129]), .D1(A[145]), .D2(A[161]), .D3(A[177]), 
        .D4(A[193]), .D5(A[209]), .D6(A[225]), .D7(A[241]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][129] ) );
    MUX81P MX8_1_5_8 ( .D0(A[136]), .D1(A[152]), .D2(A[168]), .D3(A[184]), 
        .D4(A[200]), .D5(A[216]), .D6(A[232]), .D7(A[248]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][136] ) );
    MUX81P MX8_1_5_15 ( .D0(A[143]), .D1(A[159]), .D2(A[175]), .D3(A[191]), 
        .D4(A[207]), .D5(A[223]), .D6(A[239]), .D7(A[255]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][143] ) );
    MUX81P MX8_1_5_12 ( .D0(A[140]), .D1(A[156]), .D2(A[172]), .D3(A[188]), 
        .D4(A[204]), .D5(A[220]), .D6(A[236]), .D7(A[252]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][140] ) );
    MUX81P MX8_1_1_13 ( .D0(A[13]), .D1(A[29]), .D2(A[45]), .D3(A[61]), .D4(A
        [77]), .D5(A[93]), .D6(A[109]), .D7(A[125]), .A(SEL[0]), .B(SEL[1]), 
        .C(SEL[2]), .Z(\tmp[3][13] ) );
    MUX81P MX8_1_5_6 ( .D0(A[134]), .D1(A[150]), .D2(A[166]), .D3(A[182]), 
        .D4(A[198]), .D5(A[214]), .D6(A[230]), .D7(A[246]), .A(SEL[0]), .B(SEL
        [1]), .C(SEL[2]), .Z(\tmp[3][134] ) );
    AO2 U39 ( .A(\tmp[3][9] ), .B(n58), .C(\tmp[3][137] ), .D(SEL[3]), .Z(n56)
         );
    AO2 U40 ( .A(\tmp[3][8] ), .B(n58), .C(\tmp[3][136] ), .D(SEL[3]), .Z(n59)
         );
    AO2 U41 ( .A(\tmp[3][7] ), .B(n58), .C(\tmp[3][135] ), .D(SEL[3]), .Z(n60)
         );
    AO2 U42 ( .A(\tmp[3][6] ), .B(n58), .C(\tmp[3][134] ), .D(SEL[3]), .Z(n61)
         );
    AO2 U43 ( .A(\tmp[3][5] ), .B(n58), .C(\tmp[3][133] ), .D(SEL[3]), .Z(n62)
         );
    AO2 U44 ( .A(\tmp[3][4] ), .B(n58), .C(\tmp[3][132] ), .D(SEL[3]), .Z(n63)
         );
    AO2 U45 ( .A(\tmp[3][3] ), .B(n58), .C(\tmp[3][131] ), .D(SEL[3]), .Z(n64)
         );
    AO2 U46 ( .A(\tmp[3][2] ), .B(n58), .C(\tmp[3][130] ), .D(SEL[3]), .Z(n65)
         );
    AO2 U47 ( .A(\tmp[3][1] ), .B(n58), .C(\tmp[3][129] ), .D(SEL[3]), .Z(n66)
         );
    AO2 U48 ( .A(\tmp[3][15] ), .B(n58), .C(\tmp[3][143] ), .D(SEL[3]), .Z(n67
        ) );
    AO2 U49 ( .A(\tmp[3][14] ), .B(n58), .C(\tmp[3][142] ), .D(SEL[3]), .Z(n68
        ) );
    AO2 U50 ( .A(\tmp[3][13] ), .B(n58), .C(\tmp[3][141] ), .D(SEL[3]), .Z(n69
        ) );
    AO2 U51 ( .A(\tmp[3][12] ), .B(n58), .C(\tmp[3][140] ), .D(SEL[3]), .Z(n70
        ) );
    AO2 U52 ( .A(\tmp[3][11] ), .B(n58), .C(\tmp[3][139] ), .D(SEL[3]), .Z(n71
        ) );
    AO2 U53 ( .A(\tmp[3][10] ), .B(n58), .C(\tmp[3][138] ), .D(SEL[3]), .Z(n72
        ) );
    AO2 U54 ( .A(\tmp[3][0] ), .B(n58), .C(\tmp[3][128] ), .D(SEL[3]), .Z(n73)
         );
    IV U55 ( .A(SEL[3]), .Z(n58) );
    IV U56 ( .A(n56), .Z(MUX[9]) );
    IV U57 ( .A(n59), .Z(MUX[8]) );
    IV U58 ( .A(n60), .Z(MUX[7]) );
    IV U59 ( .A(n61), .Z(MUX[6]) );
    IV U60 ( .A(n62), .Z(MUX[5]) );
    IV U61 ( .A(n63), .Z(MUX[4]) );
    IV U62 ( .A(n64), .Z(MUX[3]) );
    IV U63 ( .A(n65), .Z(MUX[2]) );
    IV U64 ( .A(n66), .Z(MUX[1]) );
    IV U65 ( .A(n67), .Z(MUX[15]) );
    IV U66 ( .A(n68), .Z(MUX[14]) );
    IV U67 ( .A(n69), .Z(MUX[13]) );
    IV U68 ( .A(n70), .Z(MUX[12]) );
    IV U69 ( .A(n71), .Z(MUX[11]) );
    IV U70 ( .A(n72), .Z(MUX[10]) );
    IV U71 ( .A(n73), .Z(MUX[0]) );
endmodule


module fifo_DW_MEM_R_W_S_LAT_16_16_0 ( clk, wr_n, rd_addr, wr_addr, data_in, 
    data_out );
output [15:0] data_out;
input  [3:0] rd_addr;
input  [15:0] wr_addr;
input  [15:0] data_in;
input  clk, wr_n;
    wire \q[15][15] , \q[15][14] , \q[15][12] , \q[15][9] , \q[15][6] , 
        \q[15][2] , \q[14][1] , \q[10][15] , \q[6][0] , \q[1][12] , 
        \din[15][0] , \q[11][13] , \q[11][9] , \q[10][3] , \din[11][2] , 
        \din[5][1] , \din[1][3] , \q[2][2] , \din[6][12] , \q[9][14] , 
        \q[8][4] , \din[0][9] , \din[10][8] , \q[6][10] , \q[3][8] , \q[3][1] , 
        \din[10][10] , \din[8][10] , \q[0][14] , \q[11][0] , \din[10][1] , 
        \din[14][3] , \din[0][0] , \din[4][2] , \q[14][8] , \q[7][3] , 
        \din[7][14] , \din[1][10] , \q[14][5] , \q[10][7] , \q[9][10] , 
        \q[9][7] , \q[8][12] , \q[6][9] , \din[15][9] , \din[5][8] , \q[8][0] , 
        \din[10][14] , \din[8][14] , \q[2][6] , \din[11][6] , \din[0][12] , 
        \din[15][4] , \din[1][7] , \din[5][5] , \q[10][11] , \q[7][12] , 
        \q[9][3] , \q[6][4] , \din[9][12] , \q[7][7] , \din[11][12] , 
        \din[14][7] , \din[7][10] , \din[1][14] , \q[15][4] , \q[11][4] , 
        \q[8][9] , \din[10][5] , \din[4][6] , \din[0][4] , \q[7][5] , 
        \q[6][14] , \q[3][5] , \q[0][10] , \din[14][5] , \din[7][12] , 
        \din[4][4] , \q[15][0] , \q[14][7] , \q[11][15] , \q[11][6] , 
        \din[10][7] , \q[3][7] , \din[0][6] , \q[0][12] , \q[10][5] , 
        \q[9][8] , \q[9][1] , \q[8][14] , \din[11][10] , \din[9][10] , 
        \q[2][4] , \din[6][14] , \din[0][10] , \din[11][4] , \din[1][5] , 
        \din[15][6] , \q[11][11] , \q[10][13] , \q[6][6] , \din[5][7] , 
        \q[10][8] , \q[9][12] , \q[8][2] , \q[7][10] , \q[1][14] , \q[8][10] , 
        \q[2][9] , \din[11][14] , \din[9][14] , \q[9][5] , \din[1][8] , 
        \q[3][3] , \din[11][9] , \q[11][2] , \q[6][12] , \din[10][3] , 
        \din[0][2] , \din[14][1] , \q[8][6] , \q[7][1] , \din[4][0] , 
        \din[1][12] , \q[7][8] , \din[10][12] , \q[14][3] , \q[7][14] , 
        \q[1][10] , \din[14][8] , \din[8][12] , \din[4][9] , \q[6][2] , 
        \din[15][2] , \din[5][3] , \q[12][7] , \q[10][1] , \din[11][0] , 
        \q[4][4] , \q[2][0] , \din[1][1] , \wren[8] , \din[6][10] , 
        \din[0][14] , \din[5][11] , \din[3][15] , \din[7][5] , \q[0][6] , 
        \din[13][6] , \din[3][7] , \q[14][14] , \q[13][4] , \q[4][15] , 
        \q[2][11] , \q[1][5] , \din[13][13] , \din[9][1] , \din[2][13] , 
        \din[9][8] , \din[2][4] , \q[12][10] , \q[5][13] , \din[12][5] , 
        \din[6][6] , \q[14][12] , \q[14][10] , \q[13][12] , \q[13][9] , 
        \q[5][7] , \q[1][8] , \wren[1] , \din[14][11] , \din[12][15] , 
        \din[15][13] , \din[8][2] , \din[12][8] , \din[9][5] , \q[4][11] , 
        \q[2][15] , \din[2][9] , \q[12][3] , \q[0][2] , \din[3][3] , \q[4][9] , 
        \q[4][0] , \din[13][2] , \din[7][1] , \din[8][6] , \din[5][15] , 
        \din[3][11] , \wren[5] , \din[14][15] , \din[12][11] , \din[7][8] , 
        \q[13][0] , \q[12][14] , \q[5][3] , \q[3][13] , \din[6][2] , 
        \q[5][15] , \q[1][1] , \wren[13] , \din[2][0] , \din[12][1] , 
        \din[4][13] , \q[3][11] , \q[13][10] , \q[13][2] , \q[5][1] , 
        \wren[11] , \din[6][0] , \din[2][2] , \q[12][8] , \q[1][3] , 
        \din[12][3] , \din[4][11] , \din[2][15] , \din[13][9] , \q[0][9] , 
        \din[3][8] , \q[0][0] , \wren[7] , \din[12][13] , \din[8][4] , 
        \q[15][11] , \q[15][10] , \q[13][6] , \q[12][1] , \q[4][13] , 
        \q[5][8] , \q[4][2] , \din[13][0] , \din[3][1] , \din[7][3] , 
        \din[3][13] , \din[6][9] , \q[1][7] , \wren[3] , \din[15][11] , 
        \din[9][7] , \din[13][15] , \din[14][13] , \din[8][0] , \din[4][15] , 
        \din[2][11] , \q[12][12] , \wren[15] , \din[2][6] , \din[12][7] , 
        \din[6][4] , \q[12][5] , \q[5][11] , \q[3][15] , \q[5][5] , \q[4][6] , 
        \din[15][15] , \din[13][11] , \din[9][3] , \din[7][7] , \din[5][13] , 
        \din[3][5] , \q[2][13] , \din[13][4] , \q[13][15] , \q[13][14] , 
        \q[13][7] , \q[0][4] , \wren[14] , \wren[2] , \din[8][9] , 
        \din[14][12] , \din[8][1] , \q[12][13] , \q[1][6] , \din[12][6] , 
        \din[2][7] , \din[4][14] , \din[2][10] , \q[5][10] , \q[5][4] , 
        \q[3][14] , \q[4][7] , \din[15][14] , \din[6][5] , \din[13][10] , 
        \din[9][2] , \din[7][6] , \din[5][12] , \q[2][12] , \q[0][5] , 
        \din[8][8] , \q[14][13] , \q[12][4] , \din[3][4] , \q[5][14] , 
        \q[3][10] , \din[13][5] , \din[6][1] , \q[13][3] , \q[5][0] , 
        \q[1][2] , \din[4][10] , \din[2][14] , \din[2][3] , \q[12][9] , 
        \q[0][8] , \wren[10] , \din[12][2] , \din[8][5] , \din[13][8] , 
        \q[12][0] , \wren[6] , \din[12][12] , \din[3][9] , \din[13][1] , 
        \din[3][0] , \q[15][13] , \q[14][11] , \q[13][13] , \q[13][11] , 
        \q[13][8] , \q[5][9] , \q[4][12] , \q[4][3] , \q[0][1] , \din[7][2] , 
        \din[3][12] , \din[15][10] , \din[13][14] , \din[9][6] , \din[6][8] , 
        \din[12][9] , \q[12][2] , \q[1][9] , \din[15][12] , \din[2][8] , 
        \din[9][4] , \din[3][2] , \q[4][10] , \q[0][3] , \din[13][3] , 
        \q[2][14] , \q[12][15] , \q[4][8] , \q[4][1] , \din[5][14] , 
        \din[3][10] , \din[8][7] , \din[7][0] , \din[7][9] , \wren[4] , 
        \din[14][14] , \din[12][10] , \din[6][3] , \q[13][1] , \q[5][2] , 
        \q[3][12] , \q[1][0] , \din[4][12] , \wren[12] , \q[4][5] , \wren[9] , 
        \din[12][0] , \din[2][1] , \din[7][4] , \din[5][10] , \din[3][14] , 
        \q[15][8] , \q[15][1] , \q[14][15] , \q[13][5] , \q[12][6] , 
        \q[4][14] , \q[2][10] , \q[0][7] , \din[13][12] , \din[13][7] , 
        \din[3][6] , \din[9][0] , \din[2][5] , \q[5][12] , \q[1][4] , 
        \din[12][4] , \din[9][9] , \din[2][12] , \q[12][11] , \q[11][10] , 
        \q[11][3] , \q[10][9] , \q[8][11] , \q[5][6] , \din[6][7] , \wren[0] , 
        \din[14][10] , \din[12][14] , \din[8][3] , \q[9][4] , \din[9][15] , 
        \q[2][8] , \din[11][15] , \din[11][8] , \din[1][9] , \din[10][2] , 
        \din[0][3] , \q[3][2] , \q[7][0] , \q[6][13] , \din[14][0] , 
        \din[1][13] , \q[8][7] , \din[4][1] , \q[15][7] , \q[15][5] , 
        \q[14][2] , \q[7][9] , \din[14][9] , \din[8][13] , \din[4][8] , 
        \din[10][13] , \din[15][3] , \din[5][2] , \q[10][0] , \q[7][15] , 
        \q[6][3] , \q[2][1] , \q[1][11] , \din[6][11] , \din[0][15] , 
        \din[11][1] , \din[14][4] , \din[1][0] , \din[4][5] , \q[14][6] , 
        \q[11][14] , \q[7][4] , \q[3][6] , \din[7][13] , \q[0][13] , 
        \q[11][7] , \din[10][6] , \q[10][12] , \q[10][4] , \q[9][9] , 
        \q[9][0] , \din[11][11] , \din[0][7] , \q[8][15] , \din[9][11] , 
        \din[11][5] , \din[1][4] , \q[2][5] , \din[6][15] , \din[0][11] , 
        \q[7][11] , \q[1][15] , \q[6][7] , \din[15][7] , \q[14][4] , 
        \q[10][10] , \q[10][6] , \q[9][13] , \q[8][3] , \din[5][6] , 
        \q[9][11] , \q[8][1] , \din[10][15] , \din[8][15] , \din[11][7] , 
        \q[7][13] , \q[6][5] , \q[2][7] , \din[1][6] , \din[0][13] , 
        \din[15][5] , \din[5][4] , \q[9][2] , \din[11][13] , \din[9][13] , 
        \din[14][6] , \q[15][3] , \q[14][0] , \q[11][5] , \q[8][8] , \q[7][6] , 
        \din[4][7] , \q[6][15] , \q[3][4] , \din[7][11] , \din[1][15] , 
        \q[0][11] , \din[10][4] , \din[0][5] , \din[15][1] , \q[11][12] , 
        \q[11][8] , \q[10][14] , \din[5][0] , \q[10][2] , \q[6][1] , 
        \q[1][13] , \q[2][3] , \din[11][3] , \din[6][13] , \din[1][2] , 
        \q[3][9] , \q[11][1] , \q[9][15] , \q[8][5] , \din[0][8] , 
        \din[10][11] , \din[10][9] , \din[8][11] , \din[10][0] , \q[6][11] , 
        \q[3][0] , \din[0][1] , \q[0][15] , \q[7][2] , \din[14][2] , 
        \din[7][15] , \din[1][11] , \din[4][3] , \q[14][9] , \q[6][8] , 
        \q[9][6] , \q[8][13] , \din[15][8] , \din[5][9] , n73, n74, n75, n76, 
        n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89;
    fifo_DW01_mux_any_256_4_16_0 MX ( .A({\q[15][15] , \q[15][14] , 
        \q[15][13] , \q[15][12] , \q[15][11] , \q[15][10] , \q[15][9] , 
        \q[15][8] , \q[15][7] , \q[15][6] , \q[15][5] , \q[15][4] , \q[15][3] , 
        \q[15][2] , \q[15][1] , \q[15][0] , \q[14][15] , \q[14][14] , 
        \q[14][13] , \q[14][12] , \q[14][11] , \q[14][10] , \q[14][9] , 
        \q[14][8] , \q[14][7] , \q[14][6] , \q[14][5] , \q[14][4] , \q[14][3] , 
        \q[14][2] , \q[14][1] , \q[14][0] , \q[13][15] , \q[13][14] , 
        \q[13][13] , \q[13][12] , \q[13][11] , \q[13][10] , \q[13][9] , 
        \q[13][8] , \q[13][7] , \q[13][6] , \q[13][5] , \q[13][4] , \q[13][3] , 
        \q[13][2] , \q[13][1] , \q[13][0] , \q[12][15] , \q[12][14] , 
        \q[12][13] , \q[12][12] , \q[12][11] , \q[12][10] , \q[12][9] , 
        \q[12][8] , \q[12][7] , \q[12][6] , \q[12][5] , \q[12][4] , \q[12][3] , 
        \q[12][2] , \q[12][1] , \q[12][0] , \q[11][15] , \q[11][14] , 
        \q[11][13] , \q[11][12] , \q[11][11] , \q[11][10] , \q[11][9] , 
        \q[11][8] , \q[11][7] , \q[11][6] , \q[11][5] , \q[11][4] , \q[11][3] , 
        \q[11][2] , \q[11][1] , \q[11][0] , \q[10][15] , \q[10][14] , 
        \q[10][13] , \q[10][12] , \q[10][11] , \q[10][10] , \q[10][9] , 
        \q[10][8] , \q[10][7] , \q[10][6] , \q[10][5] , \q[10][4] , \q[10][3] , 
        \q[10][2] , \q[10][1] , \q[10][0] , \q[9][15] , \q[9][14] , \q[9][13] , 
        \q[9][12] , \q[9][11] , \q[9][10] , \q[9][9] , \q[9][8] , \q[9][7] , 
        \q[9][6] , \q[9][5] , \q[9][4] , \q[9][3] , \q[9][2] , \q[9][1] , 
        \q[9][0] , \q[8][15] , \q[8][14] , \q[8][13] , \q[8][12] , \q[8][11] , 
        \q[8][10] , \q[8][9] , \q[8][8] , \q[8][7] , \q[8][6] , \q[8][5] , 
        \q[8][4] , \q[8][3] , \q[8][2] , \q[8][1] , \q[8][0] , \q[7][15] , 
        \q[7][14] , \q[7][13] , \q[7][12] , \q[7][11] , \q[7][10] , \q[7][9] , 
        \q[7][8] , \q[7][7] , \q[7][6] , \q[7][5] , \q[7][4] , \q[7][3] , 
        \q[7][2] , \q[7][1] , \q[7][0] , \q[6][15] , \q[6][14] , \q[6][13] , 
        \q[6][12] , \q[6][11] , \q[6][10] , \q[6][9] , \q[6][8] , \q[6][7] , 
        \q[6][6] , \q[6][5] , \q[6][4] , \q[6][3] , \q[6][2] , \q[6][1] , 
        \q[6][0] , \q[5][15] , \q[5][14] , \q[5][13] , \q[5][12] , \q[5][11] , 
        \q[5][10] , \q[5][9] , \q[5][8] , \q[5][7] , \q[5][6] , \q[5][5] , 
        \q[5][4] , \q[5][3] , \q[5][2] , \q[5][1] , \q[5][0] , \q[4][15] , 
        \q[4][14] , \q[4][13] , \q[4][12] , \q[4][11] , \q[4][10] , \q[4][9] , 
        \q[4][8] , \q[4][7] , \q[4][6] , \q[4][5] , \q[4][4] , \q[4][3] , 
        \q[4][2] , \q[4][1] , \q[4][0] , \q[3][15] , \q[3][14] , \q[3][13] , 
        \q[3][12] , \q[3][11] , \q[3][10] , \q[3][9] , \q[3][8] , \q[3][7] , 
        \q[3][6] , \q[3][5] , \q[3][4] , \q[3][3] , \q[3][2] , \q[3][1] , 
        \q[3][0] , \q[2][15] , \q[2][14] , \q[2][13] , \q[2][12] , \q[2][11] , 
        \q[2][10] , \q[2][9] , \q[2][8] , \q[2][7] , \q[2][6] , \q[2][5] , 
        \q[2][4] , \q[2][3] , \q[2][2] , \q[2][1] , \q[2][0] , \q[1][15] , 
        \q[1][14] , \q[1][13] , \q[1][12] , \q[1][11] , \q[1][10] , \q[1][9] , 
        \q[1][8] , \q[1][7] , \q[1][6] , \q[1][5] , \q[1][4] , \q[1][3] , 
        \q[1][2] , \q[1][1] , \q[1][0] , \q[0][15] , \q[0][14] , \q[0][13] , 
        \q[0][12] , \q[0][11] , \q[0][10] , \q[0][9] , \q[0][8] , \q[0][7] , 
        \q[0][6] , \q[0][5] , \q[0][4] , \q[0][3] , \q[0][2] , \q[0][1] , 
        \q[0][0] }), .SEL(rd_addr), .MUX(data_out) );
    MUX21H MX1_0_0 ( .A(\q[0][0] ), .B(data_in[0]), .S(\wren[0] ), .Z(
        \din[0][0] ) );
    MUX21H MX1_0_11 ( .A(\q[11][0] ), .B(data_in[0]), .S(\wren[11] ), .Z(
        \din[11][0] ) );
    MUX21H MX1_8_1 ( .A(\q[1][8] ), .B(data_in[8]), .S(\wren[1] ), .Z(
        \din[1][8] ) );
    MUX21H MX1_15_9 ( .A(\q[9][15] ), .B(data_in[15]), .S(\wren[9] ), .Z(
        \din[9][15] ) );
    MUX21H MX1_12_3 ( .A(\q[3][12] ), .B(data_in[12]), .S(\wren[3] ), .Z(
        \din[3][12] ) );
    MUX21H MX1_14_12 ( .A(\q[12][14] ), .B(data_in[14]), .S(\wren[12] ), .Z(
        \din[12][14] ) );
    MUX21H MX1_5_6 ( .A(\q[6][5] ), .B(data_in[5]), .S(\wren[6] ), .Z(
        \din[6][5] ) );
    MUX21H MX1_6_14 ( .A(\q[14][6] ), .B(data_in[6]), .S(\wren[14] ), .Z(
        \din[14][6] ) );
    MUX21H MX1_1_0 ( .A(\q[0][1] ), .B(data_in[1]), .S(\wren[0] ), .Z(
        \din[0][1] ) );
    MUX21H MX1_4_6 ( .A(\q[6][4] ), .B(data_in[4]), .S(\wren[6] ), .Z(
        \din[6][4] ) );
    MUX21H MX1_1_10 ( .A(\q[10][1] ), .B(data_in[1]), .S(\wren[10] ), .Z(
        \din[10][1] ) );
    MUX21H MX1_0_9 ( .A(\q[9][0] ), .B(data_in[0]), .S(\wren[9] ), .Z(
        \din[9][0] ) );
    MUX21H MX1_4_10 ( .A(\q[10][4] ), .B(data_in[4]), .S(\wren[10] ), .Z(
        \din[10][4] ) );
    MUX21H MX1_14_9 ( .A(\q[9][14] ), .B(data_in[14]), .S(\wren[9] ), .Z(
        \din[9][14] ) );
    MUX21H MX1_7_15 ( .A(\q[15][7] ), .B(data_in[7]), .S(\wren[15] ), .Z(
        \din[15][7] ) );
    MUX21H MX1_15_13 ( .A(\q[13][15] ), .B(data_in[15]), .S(\wren[13] ), .Z(
        \din[13][15] ) );
    MUX21H MX1_9_1 ( .A(\q[1][9] ), .B(data_in[9]), .S(\wren[1] ), .Z(
        \din[1][9] ) );
    MUX21H MX1_8_8 ( .A(\q[8][8] ), .B(data_in[8]), .S(\wren[8] ), .Z(
        \din[8][8] ) );
    MUX21H MX1_13_3 ( .A(\q[3][13] ), .B(data_in[13]), .S(\wren[3] ), .Z(
        \din[3][13] ) );
    MUX21H MX1_15_0 ( .A(\q[0][15] ), .B(data_in[15]), .S(\wren[0] ), .Z(
        \din[0][15] ) );
    MUX21H MX1_10_6 ( .A(\q[6][10] ), .B(data_in[10]), .S(\wren[6] ), .Z(
        \din[6][10] ) );
    MUX21H MX1_1_9 ( .A(\q[9][1] ), .B(data_in[1]), .S(\wren[9] ), .Z(
        \din[9][1] ) );
    MUX21H MX1_2_5 ( .A(\q[5][2] ), .B(data_in[2]), .S(\wren[5] ), .Z(
        \din[5][2] ) );
    MUX21H MX1_8_13 ( .A(\q[13][8] ), .B(data_in[8]), .S(\wren[13] ), .Z(
        \din[13][8] ) );
    MUX21H MX1_2_15 ( .A(\q[15][2] ), .B(data_in[2]), .S(\wren[15] ), .Z(
        \din[15][2] ) );
    MUX21H MX1_7_3 ( .A(\q[3][7] ), .B(data_in[7]), .S(\wren[3] ), .Z(
        \din[3][7] ) );
    MUX21H MX1_10_13 ( .A(\q[13][10] ), .B(data_in[10]), .S(\wren[13] ), .Z(
        \din[13][10] ) );
    MUX21H MX1_5_11 ( .A(\q[11][5] ), .B(data_in[5]), .S(\wren[11] ), .Z(
        \din[11][5] ) );
    MUX21H MX1_6_3 ( .A(\q[3][6] ), .B(data_in[6]), .S(\wren[3] ), .Z(
        \din[3][6] ) );
    MUX21H MX1_3_5 ( .A(\q[5][3] ), .B(data_in[3]), .S(\wren[5] ), .Z(
        \din[5][3] ) );
    MUX21H MX1_3_14 ( .A(\q[14][3] ), .B(data_in[3]), .S(\wren[14] ), .Z(
        \din[14][3] ) );
    MUX21H MX1_9_8 ( .A(\q[8][9] ), .B(data_in[9]), .S(\wren[8] ), .Z(
        \din[8][9] ) );
    MUX21H MX1_9_12 ( .A(\q[12][9] ), .B(data_in[9]), .S(\wren[12] ), .Z(
        \din[12][9] ) );
    MUX21H MX1_11_6 ( .A(\q[6][11] ), .B(data_in[11]), .S(\wren[6] ), .Z(
        \din[6][11] ) );
    MUX21H MX1_14_0 ( .A(\q[0][14] ), .B(data_in[14]), .S(\wren[0] ), .Z(
        \din[0][14] ) );
    MUX21H MX1_9_15 ( .A(\q[15][9] ), .B(data_in[9]), .S(\wren[15] ), .Z(
        \din[15][9] ) );
    MUX21H MX1_11_12 ( .A(\q[12][11] ), .B(data_in[11]), .S(\wren[12] ), .Z(
        \din[12][11] ) );
    MUX21H MX1_14_7 ( .A(\q[7][14] ), .B(data_in[14]), .S(\wren[7] ), .Z(
        \din[7][14] ) );
    MUX21H MX1_11_1 ( .A(\q[1][11] ), .B(data_in[11]), .S(\wren[1] ), .Z(
        \din[1][11] ) );
    MUX21H MX1_3_13 ( .A(\q[13][3] ), .B(data_in[3]), .S(\wren[13] ), .Z(
        \din[13][3] ) );
    MUX21H MX1_11_15 ( .A(\q[15][11] ), .B(data_in[11]), .S(\wren[15] ), .Z(
        \din[15][11] ) );
    MUX21H MX1_4_8 ( .A(\q[8][4] ), .B(data_in[4]), .S(\wren[8] ), .Z(
        \din[8][4] ) );
    MUX21H MX1_3_2 ( .A(\q[2][3] ), .B(data_in[3]), .S(\wren[2] ), .Z(
        \din[2][3] ) );
    MUX21H MX1_6_4 ( .A(\q[4][6] ), .B(data_in[6]), .S(\wren[4] ), .Z(
        \din[4][6] ) );
    MUX21H MX1_2_2 ( .A(\q[2][2] ), .B(data_in[2]), .S(\wren[2] ), .Z(
        \din[2][2] ) );
    MUX21H MX1_2_12 ( .A(\q[12][2] ), .B(data_in[2]), .S(\wren[12] ), .Z(
        \din[12][2] ) );
    MUX21H MX1_5_8 ( .A(\q[8][5] ), .B(data_in[5]), .S(\wren[8] ), .Z(
        \din[8][5] ) );
    MUX21H MX1_8_14 ( .A(\q[14][8] ), .B(data_in[8]), .S(\wren[14] ), .Z(
        \din[14][8] ) );
    MUX21H MX1_10_14 ( .A(\q[14][10] ), .B(data_in[10]), .S(\wren[14] ), .Z(
        \din[14][10] ) );
    MUX21H MX1_7_4 ( .A(\q[4][7] ), .B(data_in[7]), .S(\wren[4] ), .Z(
        \din[4][7] ) );
    MUX21H MX1_7_12 ( .A(\q[12][7] ), .B(data_in[7]), .S(\wren[12] ), .Z(
        \din[12][7] ) );
    MUX21H MX1_10_1 ( .A(\q[1][10] ), .B(data_in[10]), .S(\wren[1] ), .Z(
        \din[1][10] ) );
    MUX21H MX1_15_7 ( .A(\q[7][15] ), .B(data_in[15]), .S(\wren[7] ), .Z(
        \din[7][15] ) );
    MUX21H MX1_9_6 ( .A(\q[6][9] ), .B(data_in[9]), .S(\wren[6] ), .Z(
        \din[6][9] ) );
    MUX21H MX1_11_8 ( .A(\q[8][11] ), .B(data_in[11]), .S(\wren[8] ), .Z(
        \din[8][11] ) );
    MUX21H MX1_13_4 ( .A(\q[4][13] ), .B(data_in[13]), .S(\wren[4] ), .Z(
        \din[4][13] ) );
    MUX21H MX1_15_14 ( .A(\q[14][15] ), .B(data_in[15]), .S(\wren[14] ), .Z(
        \din[14][15] ) );
    MUX21H MX1_0_1 ( .A(\q[1][0] ), .B(data_in[0]), .S(\wren[1] ), .Z(
        \din[1][0] ) );
    MUX21H MX1_0_6 ( .A(\q[6][0] ), .B(data_in[0]), .S(\wren[6] ), .Z(
        \din[6][0] ) );
    MUX21H MX1_0_7 ( .A(\q[7][0] ), .B(data_in[0]), .S(\wren[7] ), .Z(
        \din[7][0] ) );
    MUX21H MX1_1_7 ( .A(\q[7][1] ), .B(data_in[1]), .S(\wren[7] ), .Z(
        \din[7][1] ) );
    MUX21H MX1_4_1 ( .A(\q[1][4] ), .B(data_in[4]), .S(\wren[1] ), .Z(
        \din[1][4] ) );
    MUX21H MX1_13_11 ( .A(\q[11][13] ), .B(data_in[13]), .S(\wren[11] ), .Z(
        \din[11][13] ) );
    MUX21H MX1_5_1 ( .A(\q[1][5] ), .B(data_in[5]), .S(\wren[1] ), .Z(
        \din[1][5] ) );
    MUX21H MX1_6_13 ( .A(\q[13][6] ), .B(data_in[6]), .S(\wren[13] ), .Z(
        \din[13][6] ) );
    MUX21H MX1_14_15 ( .A(\q[15][14] ), .B(data_in[14]), .S(\wren[15] ), .Z(
        \din[15][14] ) );
    MUX21H MX1_8_6 ( .A(\q[6][8] ), .B(data_in[8]), .S(\wren[6] ), .Z(
        \din[6][8] ) );
    MUX21H MX1_8_15 ( .A(\q[15][8] ), .B(data_in[8]), .S(\wren[15] ), .Z(
        \din[15][8] ) );
    MUX21H MX1_10_8 ( .A(\q[8][10] ), .B(data_in[10]), .S(\wren[8] ), .Z(
        \din[8][10] ) );
    MUX21H MX1_12_10 ( .A(\q[10][12] ), .B(data_in[12]), .S(\wren[10] ), .Z(
        \din[10][12] ) );
    MUX21H MX1_12_4 ( .A(\q[4][12] ), .B(data_in[12]), .S(\wren[4] ), .Z(
        \din[4][12] ) );
    MUX21H MX1_10_0 ( .A(\q[0][10] ), .B(data_in[10]), .S(\wren[0] ), .Z(
        \din[0][10] ) );
    MUX21H MX1_15_6 ( .A(\q[6][15] ), .B(data_in[15]), .S(\wren[6] ), .Z(
        \din[6][15] ) );
    MUX21H MX1_2_3 ( .A(\q[3][2] ), .B(data_in[2]), .S(\wren[3] ), .Z(
        \din[3][2] ) );
    MUX21H MX1_2_13 ( .A(\q[13][2] ), .B(data_in[2]), .S(\wren[13] ), .Z(
        \din[13][2] ) );
    MUX21H MX1_5_9 ( .A(\q[9][5] ), .B(data_in[5]), .S(\wren[9] ), .Z(
        \din[9][5] ) );
    MUX21H MX1_7_5 ( .A(\q[5][7] ), .B(data_in[7]), .S(\wren[5] ), .Z(
        \din[5][7] ) );
    MUX21H MX1_10_15 ( .A(\q[15][10] ), .B(data_in[10]), .S(\wren[15] ), .Z(
        \din[15][10] ) );
    MUX21H MX1_4_9 ( .A(\q[9][4] ), .B(data_in[4]), .S(\wren[9] ), .Z(
        \din[9][4] ) );
    MUX21H MX1_3_3 ( .A(\q[3][3] ), .B(data_in[3]), .S(\wren[3] ), .Z(
        \din[3][3] ) );
    MUX21H MX1_6_5 ( .A(\q[5][6] ), .B(data_in[6]), .S(\wren[5] ), .Z(
        \din[5][6] ) );
    MUX21H MX1_9_14 ( .A(\q[14][9] ), .B(data_in[9]), .S(\wren[14] ), .Z(
        \din[14][9] ) );
    MUX21H MX1_14_6 ( .A(\q[6][14] ), .B(data_in[14]), .S(\wren[6] ), .Z(
        \din[6][14] ) );
    MUX21H MX1_11_0 ( .A(\q[0][11] ), .B(data_in[11]), .S(\wren[0] ), .Z(
        \din[0][11] ) );
    MUX21H MX1_3_12 ( .A(\q[12][3] ), .B(data_in[3]), .S(\wren[12] ), .Z(
        \din[12][3] ) );
    MUX21H MX1_11_14 ( .A(\q[14][11] ), .B(data_in[11]), .S(\wren[14] ), .Z(
        \din[14][11] ) );
    MUX21H MX1_5_0 ( .A(\q[0][5] ), .B(data_in[5]), .S(\wren[0] ), .Z(
        \din[0][5] ) );
    MUX21H MX1_8_7 ( .A(\q[7][8] ), .B(data_in[8]), .S(\wren[7] ), .Z(
        \din[7][8] ) );
    MUX21H MX1_10_9 ( .A(\q[9][10] ), .B(data_in[10]), .S(\wren[9] ), .Z(
        \din[9][10] ) );
    MUX21H MX1_12_11 ( .A(\q[11][12] ), .B(data_in[12]), .S(\wren[11] ), .Z(
        \din[11][12] ) );
    MUX21H MX1_12_5 ( .A(\q[5][12] ), .B(data_in[12]), .S(\wren[5] ), .Z(
        \din[5][12] ) );
    MUX21H MX1_6_12 ( .A(\q[12][6] ), .B(data_in[6]), .S(\wren[12] ), .Z(
        \din[12][6] ) );
    MUX21H MX1_14_14 ( .A(\q[14][14] ), .B(data_in[14]), .S(\wren[14] ), .Z(
        \din[14][14] ) );
    MUX21H MX1_1_6 ( .A(\q[6][1] ), .B(data_in[1]), .S(\wren[6] ), .Z(
        \din[6][1] ) );
    MUX21H MX1_4_0 ( .A(\q[0][4] ), .B(data_in[4]), .S(\wren[0] ), .Z(
        \din[0][4] ) );
    MUX21H MX1_7_13 ( .A(\q[13][7] ), .B(data_in[7]), .S(\wren[13] ), .Z(
        \din[13][7] ) );
    MUX21H MX1_13_10 ( .A(\q[10][13] ), .B(data_in[13]), .S(\wren[10] ), .Z(
        \din[10][13] ) );
    MUX21H MX1_11_9 ( .A(\q[9][11] ), .B(data_in[11]), .S(\wren[9] ), .Z(
        \din[9][11] ) );
    MUX21H MX1_9_7 ( .A(\q[7][9] ), .B(data_in[9]), .S(\wren[7] ), .Z(
        \din[7][9] ) );
    MUX21H MX1_13_5 ( .A(\q[5][13] ), .B(data_in[13]), .S(\wren[5] ), .Z(
        \din[5][13] ) );
    MUX21H MX1_15_15 ( .A(\q[15][15] ), .B(data_in[15]), .S(\wren[15] ), .Z(
        \din[15][15] ) );
    MUX21H MX1_7_14 ( .A(\q[14][7] ), .B(data_in[7]), .S(\wren[14] ), .Z(
        \din[14][7] ) );
    MUX21H MX1_9_0 ( .A(\q[0][9] ), .B(data_in[9]), .S(\wren[0] ), .Z(
        \din[0][9] ) );
    MUX21H MX1_14_8 ( .A(\q[8][14] ), .B(data_in[14]), .S(\wren[8] ), .Z(
        \din[8][14] ) );
    MUX21H MX1_15_12 ( .A(\q[12][15] ), .B(data_in[15]), .S(\wren[12] ), .Z(
        \din[12][15] ) );
    MUX21H MX1_13_2 ( .A(\q[2][13] ), .B(data_in[13]), .S(\wren[2] ), .Z(
        \din[2][13] ) );
    MUX21H MX1_1_1 ( .A(\q[1][1] ), .B(data_in[1]), .S(\wren[1] ), .Z(
        \din[1][1] ) );
    MUX21H MX1_1_11 ( .A(\q[11][1] ), .B(data_in[1]), .S(\wren[11] ), .Z(
        \din[11][1] ) );
    MUX21H MX1_4_7 ( .A(\q[7][4] ), .B(data_in[4]), .S(\wren[7] ), .Z(
        \din[7][4] ) );
    MUX21H MX1_14_13 ( .A(\q[13][14] ), .B(data_in[14]), .S(\wren[13] ), .Z(
        \din[13][14] ) );
    MUX21H MX1_0_2 ( .A(\q[2][0] ), .B(data_in[0]), .S(\wren[2] ), .Z(
        \din[2][0] ) );
    MUX21H MX1_0_3 ( .A(\q[3][0] ), .B(data_in[0]), .S(\wren[3] ), .Z(
        \din[3][0] ) );
    MUX21H MX1_0_8 ( .A(\q[8][0] ), .B(data_in[0]), .S(\wren[8] ), .Z(
        \din[8][0] ) );
    MUX21H MX1_0_10 ( .A(\q[10][0] ), .B(data_in[0]), .S(\wren[10] ), .Z(
        \din[10][0] ) );
    MUX21H MX1_5_7 ( .A(\q[7][5] ), .B(data_in[5]), .S(\wren[7] ), .Z(
        \din[7][5] ) );
    MUX21H MX1_6_15 ( .A(\q[15][6] ), .B(data_in[6]), .S(\wren[15] ), .Z(
        \din[15][6] ) );
    MUX21H MX1_8_0 ( .A(\q[0][8] ), .B(data_in[8]), .S(\wren[0] ), .Z(
        \din[0][8] ) );
    MUX21H MX1_1_8 ( .A(\q[8][1] ), .B(data_in[1]), .S(\wren[8] ), .Z(
        \din[8][1] ) );
    MUX21H MX1_3_15 ( .A(\q[15][3] ), .B(data_in[3]), .S(\wren[15] ), .Z(
        \din[15][3] ) );
    MUX21H MX1_12_2 ( .A(\q[2][12] ), .B(data_in[12]), .S(\wren[2] ), .Z(
        \din[2][12] ) );
    MUX21H MX1_15_8 ( .A(\q[8][15] ), .B(data_in[15]), .S(\wren[8] ), .Z(
        \din[8][15] ) );
    MUX21H MX1_9_9 ( .A(\q[9][9] ), .B(data_in[9]), .S(\wren[9] ), .Z(
        \din[9][9] ) );
    MUX21H MX1_11_7 ( .A(\q[7][11] ), .B(data_in[11]), .S(\wren[7] ), .Z(
        \din[7][11] ) );
    MUX21H MX1_9_13 ( .A(\q[13][9] ), .B(data_in[9]), .S(\wren[13] ), .Z(
        \din[13][9] ) );
    MUX21H MX1_14_1 ( .A(\q[1][14] ), .B(data_in[14]), .S(\wren[1] ), .Z(
        \din[1][14] ) );
    MUX21H MX1_11_13 ( .A(\q[13][11] ), .B(data_in[11]), .S(\wren[13] ), .Z(
        \din[13][11] ) );
    MUX21H MX1_5_10 ( .A(\q[10][5] ), .B(data_in[5]), .S(\wren[10] ), .Z(
        \din[10][5] ) );
    MUX21H MX1_6_2 ( .A(\q[2][6] ), .B(data_in[6]), .S(\wren[2] ), .Z(
        \din[2][6] ) );
    MUX21H MX1_3_4 ( .A(\q[4][3] ), .B(data_in[3]), .S(\wren[4] ), .Z(
        \din[4][3] ) );
    MUX21H MX1_0_12 ( .A(\q[12][0] ), .B(data_in[0]), .S(\wren[12] ), .Z(
        \din[12][0] ) );
    MUX21H MX1_2_4 ( .A(\q[4][2] ), .B(data_in[2]), .S(\wren[4] ), .Z(
        \din[4][2] ) );
    MUX21H MX1_8_12 ( .A(\q[12][8] ), .B(data_in[8]), .S(\wren[12] ), .Z(
        \din[12][8] ) );
    MUX21H MX1_2_14 ( .A(\q[14][2] ), .B(data_in[2]), .S(\wren[14] ), .Z(
        \din[14][2] ) );
    MUX21H MX1_7_2 ( .A(\q[2][7] ), .B(data_in[7]), .S(\wren[2] ), .Z(
        \din[2][7] ) );
    MUX21H MX1_4_11 ( .A(\q[11][4] ), .B(data_in[4]), .S(\wren[11] ), .Z(
        \din[11][4] ) );
    MUX21H MX1_10_12 ( .A(\q[12][10] ), .B(data_in[10]), .S(\wren[12] ), .Z(
        \din[12][10] ) );
    MUX21H MX1_8_9 ( .A(\q[9][8] ), .B(data_in[8]), .S(\wren[9] ), .Z(
        \din[9][8] ) );
    MUX21H MX1_10_7 ( .A(\q[7][10] ), .B(data_in[10]), .S(\wren[7] ), .Z(
        \din[7][10] ) );
    MUX21H MX1_15_1 ( .A(\q[1][15] ), .B(data_in[15]), .S(\wren[1] ), .Z(
        \din[1][15] ) );
    MUX21H MX1_12_0 ( .A(\q[0][12] ), .B(data_in[12]), .S(\wren[0] ), .Z(
        \din[0][12] ) );
    MUX21H MX1_8_2 ( .A(\q[2][8] ), .B(data_in[8]), .S(\wren[2] ), .Z(
        \din[2][8] ) );
    MUX21H MX1_12_14 ( .A(\q[14][12] ), .B(data_in[12]), .S(\wren[14] ), .Z(
        \din[14][12] ) );
    MUX21H MX1_7_9 ( .A(\q[9][7] ), .B(data_in[7]), .S(\wren[9] ), .Z(
        \din[9][7] ) );
    MUX21H MX1_5_5 ( .A(\q[5][5] ), .B(data_in[5]), .S(\wren[5] ), .Z(
        \din[5][5] ) );
    MUX21H MX1_1_3 ( .A(\q[3][1] ), .B(data_in[1]), .S(\wren[3] ), .Z(
        \din[3][1] ) );
    MUX21H MX1_6_9 ( .A(\q[9][6] ), .B(data_in[6]), .S(\wren[9] ), .Z(
        \din[9][6] ) );
    MUX21H MX1_14_11 ( .A(\q[11][14] ), .B(data_in[14]), .S(\wren[11] ), .Z(
        \din[11][14] ) );
    MUX21H MX1_1_13 ( .A(\q[13][1] ), .B(data_in[1]), .S(\wren[13] ), .Z(
        \din[13][1] ) );
    MUX21H MX1_2_1 ( .A(\q[1][2] ), .B(data_in[2]), .S(\wren[1] ), .Z(
        \din[1][2] ) );
    MUX21H MX1_2_6 ( .A(\q[6][2] ), .B(data_in[2]), .S(\wren[6] ), .Z(
        \din[6][2] ) );
    MUX21H MX1_4_5 ( .A(\q[5][4] ), .B(data_in[4]), .S(\wren[5] ), .Z(
        \din[5][4] ) );
    MUX21H MX1_13_15 ( .A(\q[15][13] ), .B(data_in[13]), .S(\wren[15] ), .Z(
        \din[15][13] ) );
    MUX21H MX1_4_13 ( .A(\q[13][4] ), .B(data_in[4]), .S(\wren[13] ), .Z(
        \din[13][4] ) );
    MUX21H MX1_9_2 ( .A(\q[2][9] ), .B(data_in[9]), .S(\wren[2] ), .Z(
        \din[2][9] ) );
    MUX21H MX1_13_0 ( .A(\q[0][13] ), .B(data_in[13]), .S(\wren[0] ), .Z(
        \din[0][13] ) );
    MUX21H MX1_15_10 ( .A(\q[10][15] ), .B(data_in[15]), .S(\wren[10] ), .Z(
        \din[10][15] ) );
    MUX21H MX1_12_9 ( .A(\q[9][12] ), .B(data_in[12]), .S(\wren[9] ), .Z(
        \din[9][12] ) );
    MUX21H MX1_7_0 ( .A(\q[0][7] ), .B(data_in[7]), .S(\wren[0] ), .Z(
        \din[0][7] ) );
    MUX21H MX1_10_5 ( .A(\q[5][10] ), .B(data_in[10]), .S(\wren[5] ), .Z(
        \din[5][10] ) );
    MUX21H MX1_15_3 ( .A(\q[3][15] ), .B(data_in[15]), .S(\wren[3] ), .Z(
        \din[3][15] ) );
    MUX21H MX1_10_10 ( .A(\q[10][10] ), .B(data_in[10]), .S(\wren[10] ), .Z(
        \din[10][10] ) );
    MUX21H MX1_8_10 ( .A(\q[10][8] ), .B(data_in[8]), .S(\wren[10] ), .Z(
        \din[10][8] ) );
    MUX21H MX1_3_6 ( .A(\q[6][3] ), .B(data_in[3]), .S(\wren[6] ), .Z(
        \din[6][3] ) );
    MUX21H MX1_3_10 ( .A(\q[10][3] ), .B(data_in[3]), .S(\wren[10] ), .Z(
        \din[10][3] ) );
    MUX21H MX1_5_12 ( .A(\q[12][5] ), .B(data_in[5]), .S(\wren[12] ), .Z(
        \din[12][5] ) );
    MUX21H MX1_6_0 ( .A(\q[0][6] ), .B(data_in[6]), .S(\wren[0] ), .Z(
        \din[0][6] ) );
    MUX21H MX1_9_11 ( .A(\q[11][9] ), .B(data_in[9]), .S(\wren[11] ), .Z(
        \din[11][9] ) );
    MUX21H MX1_11_11 ( .A(\q[11][11] ), .B(data_in[11]), .S(\wren[11] ), .Z(
        \din[11][11] ) );
    MUX21H MX1_13_9 ( .A(\q[9][13] ), .B(data_in[13]), .S(\wren[9] ), .Z(
        \din[9][13] ) );
    MUX21H MX1_14_3 ( .A(\q[3][14] ), .B(data_in[14]), .S(\wren[3] ), .Z(
        \din[3][14] ) );
    MUX21H MX1_11_5 ( .A(\q[5][11] ), .B(data_in[11]), .S(\wren[5] ), .Z(
        \din[5][11] ) );
    MUX21H MX1_3_1 ( .A(\q[1][3] ), .B(data_in[3]), .S(\wren[1] ), .Z(
        \din[1][3] ) );
    MUX21H MX1_5_15 ( .A(\q[15][5] ), .B(data_in[5]), .S(\wren[15] ), .Z(
        \din[15][5] ) );
    MUX21H MX1_6_7 ( .A(\q[7][6] ), .B(data_in[6]), .S(\wren[7] ), .Z(
        \din[7][6] ) );
    MUX21H MX1_11_2 ( .A(\q[2][11] ), .B(data_in[11]), .S(\wren[2] ), .Z(
        \din[2][11] ) );
    MUX21H MX1_14_4 ( .A(\q[4][14] ), .B(data_in[14]), .S(\wren[4] ), .Z(
        \din[4][14] ) );
    MUX21H MX1_2_11 ( .A(\q[11][2] ), .B(data_in[2]), .S(\wren[11] ), .Z(
        \din[11][2] ) );
    MUX21H MX1_3_8 ( .A(\q[8][3] ), .B(data_in[3]), .S(\wren[8] ), .Z(
        \din[8][3] ) );
    MUX21H MX1_4_14 ( .A(\q[14][4] ), .B(data_in[4]), .S(\wren[14] ), .Z(
        \din[14][4] ) );
    MUX21H MX1_7_7 ( .A(\q[7][7] ), .B(data_in[7]), .S(\wren[7] ), .Z(
        \din[7][7] ) );
    MUX21H MX1_10_2 ( .A(\q[2][10] ), .B(data_in[10]), .S(\wren[2] ), .Z(
        \din[2][10] ) );
    MUX21H MX1_15_4 ( .A(\q[4][15] ), .B(data_in[15]), .S(\wren[4] ), .Z(
        \din[4][15] ) );
    MUX21H MX1_13_7 ( .A(\q[7][13] ), .B(data_in[13]), .S(\wren[7] ), .Z(
        \din[7][13] ) );
    MUX21H MX1_7_11 ( .A(\q[11][7] ), .B(data_in[7]), .S(\wren[11] ), .Z(
        \din[11][7] ) );
    MUX21H MX1_9_5 ( .A(\q[5][9] ), .B(data_in[9]), .S(\wren[5] ), .Z(
        \din[5][9] ) );
    MUX21H MX1_4_2 ( .A(\q[2][4] ), .B(data_in[4]), .S(\wren[2] ), .Z(
        \din[2][4] ) );
    MUX21H MX1_13_12 ( .A(\q[12][13] ), .B(data_in[13]), .S(\wren[12] ), .Z(
        \din[12][13] ) );
    MUX21H MX1_0_4 ( .A(\q[4][0] ), .B(data_in[0]), .S(\wren[4] ), .Z(
        \din[4][0] ) );
    MUX21H MX1_1_4 ( .A(\q[4][1] ), .B(data_in[1]), .S(\wren[4] ), .Z(
        \din[4][1] ) );
    MUX21H MX1_1_14 ( .A(\q[14][1] ), .B(data_in[1]), .S(\wren[14] ), .Z(
        \din[14][1] ) );
    MUX21H MX1_2_8 ( .A(\q[8][2] ), .B(data_in[2]), .S(\wren[8] ), .Z(
        \din[8][2] ) );
    MUX21H MX1_0_5 ( .A(\q[5][0] ), .B(data_in[0]), .S(\wren[5] ), .Z(
        \din[5][0] ) );
    MUX21H MX1_0_14 ( .A(\q[14][0] ), .B(data_in[0]), .S(\wren[14] ), .Z(
        \din[14][0] ) );
    MUX21H MX1_0_15 ( .A(\q[15][0] ), .B(data_in[0]), .S(\wren[15] ), .Z(
        \din[15][0] ) );
    MUX21H MX1_5_2 ( .A(\q[2][5] ), .B(data_in[5]), .S(\wren[2] ), .Z(
        \din[2][5] ) );
    MUX21H MX1_6_10 ( .A(\q[10][6] ), .B(data_in[6]), .S(\wren[10] ), .Z(
        \din[10][6] ) );
    MUX21H MX1_8_5 ( .A(\q[5][8] ), .B(data_in[8]), .S(\wren[5] ), .Z(
        \din[5][8] ) );
    MUX21H MX1_12_7 ( .A(\q[7][12] ), .B(data_in[12]), .S(\wren[7] ), .Z(
        \din[7][12] ) );
    MUX21H MX1_12_13 ( .A(\q[13][12] ), .B(data_in[12]), .S(\wren[13] ), .Z(
        \din[13][12] ) );
    MUX21H MX1_2_0 ( .A(\q[0][2] ), .B(data_in[2]), .S(\wren[0] ), .Z(
        \din[0][2] ) );
    MUX21H MX1_2_10 ( .A(\q[10][2] ), .B(data_in[2]), .S(\wren[10] ), .Z(
        \din[10][2] ) );
    MUX21H MX1_4_15 ( .A(\q[15][4] ), .B(data_in[4]), .S(\wren[15] ), .Z(
        \din[15][4] ) );
    MUX21H MX1_10_3 ( .A(\q[3][10] ), .B(data_in[10]), .S(\wren[3] ), .Z(
        \din[3][10] ) );
    MUX21H MX1_15_5 ( .A(\q[5][15] ), .B(data_in[15]), .S(\wren[5] ), .Z(
        \din[5][15] ) );
    MUX21H MX1_3_0 ( .A(\q[0][3] ), .B(data_in[3]), .S(\wren[0] ), .Z(
        \din[0][3] ) );
    MUX21H MX1_5_14 ( .A(\q[14][5] ), .B(data_in[5]), .S(\wren[14] ), .Z(
        \din[14][5] ) );
    MUX21H MX1_6_6 ( .A(\q[6][6] ), .B(data_in[6]), .S(\wren[6] ), .Z(
        \din[6][6] ) );
    MUX21H MX1_7_6 ( .A(\q[6][7] ), .B(data_in[7]), .S(\wren[6] ), .Z(
        \din[6][7] ) );
    MUX21H MX1_3_11 ( .A(\q[11][3] ), .B(data_in[3]), .S(\wren[11] ), .Z(
        \din[11][3] ) );
    MUX21H MX1_11_3 ( .A(\q[3][11] ), .B(data_in[11]), .S(\wren[3] ), .Z(
        \din[3][11] ) );
    MUX21H MX1_12_6 ( .A(\q[6][12] ), .B(data_in[12]), .S(\wren[6] ), .Z(
        \din[6][12] ) );
    MUX21H MX1_14_5 ( .A(\q[5][14] ), .B(data_in[14]), .S(\wren[5] ), .Z(
        \din[5][14] ) );
    MUX21H MX1_8_4 ( .A(\q[4][8] ), .B(data_in[8]), .S(\wren[4] ), .Z(
        \din[4][8] ) );
    MUX21H MX1_12_12 ( .A(\q[12][12] ), .B(data_in[12]), .S(\wren[12] ), .Z(
        \din[12][12] ) );
    MUX21H MX1_2_9 ( .A(\q[9][2] ), .B(data_in[2]), .S(\wren[9] ), .Z(
        \din[9][2] ) );
    MUX21H MX1_3_9 ( .A(\q[9][3] ), .B(data_in[3]), .S(\wren[9] ), .Z(
        \din[9][3] ) );
    MUX21H MX1_5_3 ( .A(\q[3][5] ), .B(data_in[5]), .S(\wren[3] ), .Z(
        \din[3][5] ) );
    MUX21H MX1_6_11 ( .A(\q[11][6] ), .B(data_in[6]), .S(\wren[11] ), .Z(
        \din[11][6] ) );
    MUX21H MX1_4_3 ( .A(\q[3][4] ), .B(data_in[4]), .S(\wren[3] ), .Z(
        \din[3][4] ) );
    MUX21H MX1_13_13 ( .A(\q[13][13] ), .B(data_in[13]), .S(\wren[13] ), .Z(
        \din[13][13] ) );
    MUX21H MX1_1_2 ( .A(\q[2][1] ), .B(data_in[1]), .S(\wren[2] ), .Z(
        \din[2][1] ) );
    MUX21H MX1_1_5 ( .A(\q[5][1] ), .B(data_in[1]), .S(\wren[5] ), .Z(
        \din[5][1] ) );
    MUX21H MX1_1_12 ( .A(\q[12][1] ), .B(data_in[1]), .S(\wren[12] ), .Z(
        \din[12][1] ) );
    MUX21H MX1_1_15 ( .A(\q[15][1] ), .B(data_in[1]), .S(\wren[15] ), .Z(
        \din[15][1] ) );
    MUX21H MX1_6_8 ( .A(\q[8][6] ), .B(data_in[6]), .S(\wren[8] ), .Z(
        \din[8][6] ) );
    MUX21H MX1_13_6 ( .A(\q[6][13] ), .B(data_in[13]), .S(\wren[6] ), .Z(
        \din[6][13] ) );
    MUX21H MX1_7_10 ( .A(\q[10][7] ), .B(data_in[7]), .S(\wren[10] ), .Z(
        \din[10][7] ) );
    MUX21H MX1_9_3 ( .A(\q[3][9] ), .B(data_in[9]), .S(\wren[3] ), .Z(
        \din[3][9] ) );
    MUX21H MX1_9_4 ( .A(\q[4][9] ), .B(data_in[9]), .S(\wren[4] ), .Z(
        \din[4][9] ) );
    MUX21H MX1_13_1 ( .A(\q[1][13] ), .B(data_in[13]), .S(\wren[1] ), .Z(
        \din[1][13] ) );
    MUX21H MX1_15_11 ( .A(\q[11][15] ), .B(data_in[15]), .S(\wren[11] ), .Z(
        \din[11][15] ) );
    MUX21H MX1_4_4 ( .A(\q[4][4] ), .B(data_in[4]), .S(\wren[4] ), .Z(
        \din[4][4] ) );
    MUX21H MX1_13_14 ( .A(\q[14][13] ), .B(data_in[13]), .S(\wren[14] ), .Z(
        \din[14][13] ) );
    MUX21H MX1_7_8 ( .A(\q[8][7] ), .B(data_in[7]), .S(\wren[8] ), .Z(
        \din[8][7] ) );
    MUX21H MX1_5_4 ( .A(\q[4][5] ), .B(data_in[5]), .S(\wren[4] ), .Z(
        \din[4][5] ) );
    MUX21H MX1_14_10 ( .A(\q[10][14] ), .B(data_in[14]), .S(\wren[10] ), .Z(
        \din[10][14] ) );
    MUX21H MX1_0_13 ( .A(\q[13][0] ), .B(data_in[0]), .S(\wren[13] ), .Z(
        \din[13][0] ) );
    MUX21H MX1_12_1 ( .A(\q[1][12] ), .B(data_in[12]), .S(\wren[1] ), .Z(
        \din[1][12] ) );
    MUX21H MX1_8_3 ( .A(\q[3][8] ), .B(data_in[8]), .S(\wren[3] ), .Z(
        \din[3][8] ) );
    MUX21H MX1_9_10 ( .A(\q[10][9] ), .B(data_in[9]), .S(\wren[10] ), .Z(
        \din[10][9] ) );
    MUX21H MX1_11_10 ( .A(\q[10][11] ), .B(data_in[11]), .S(\wren[10] ), .Z(
        \din[10][11] ) );
    MUX21H MX1_12_15 ( .A(\q[15][12] ), .B(data_in[12]), .S(\wren[15] ), .Z(
        \din[15][12] ) );
    MUX21H MX1_13_8 ( .A(\q[8][13] ), .B(data_in[13]), .S(\wren[8] ), .Z(
        \din[8][13] ) );
    MUX21H MX1_14_2 ( .A(\q[2][14] ), .B(data_in[14]), .S(\wren[2] ), .Z(
        \din[2][14] ) );
    MUX21H MX1_11_4 ( .A(\q[4][11] ), .B(data_in[11]), .S(\wren[4] ), .Z(
        \din[4][11] ) );
    MUX21H MX1_2_7 ( .A(\q[7][2] ), .B(data_in[2]), .S(\wren[7] ), .Z(
        \din[7][2] ) );
    MUX21H MX1_3_7 ( .A(\q[7][3] ), .B(data_in[3]), .S(\wren[7] ), .Z(
        \din[7][3] ) );
    MUX21H MX1_5_13 ( .A(\q[13][5] ), .B(data_in[5]), .S(\wren[13] ), .Z(
        \din[13][5] ) );
    MUX21H MX1_6_1 ( .A(\q[1][6] ), .B(data_in[6]), .S(\wren[1] ), .Z(
        \din[1][6] ) );
    MUX21H MX1_7_1 ( .A(\q[1][7] ), .B(data_in[7]), .S(\wren[1] ), .Z(
        \din[1][7] ) );
    MUX21H MX1_10_11 ( .A(\q[11][10] ), .B(data_in[10]), .S(\wren[11] ), .Z(
        \din[11][10] ) );
    MUX21H MX1_4_12 ( .A(\q[12][4] ), .B(data_in[4]), .S(\wren[12] ), .Z(
        \din[12][4] ) );
    MUX21H MX1_8_11 ( .A(\q[11][8] ), .B(data_in[8]), .S(\wren[11] ), .Z(
        \din[11][8] ) );
    MUX21H MX1_12_8 ( .A(\q[8][12] ), .B(data_in[12]), .S(\wren[8] ), .Z(
        \din[8][12] ) );
    MUX21H MX1_10_4 ( .A(\q[4][10] ), .B(data_in[10]), .S(\wren[4] ), .Z(
        \din[4][10] ) );
    MUX21H MX1_15_2 ( .A(\q[2][15] ), .B(data_in[15]), .S(\wren[2] ), .Z(
        \din[2][15] ) );
    LD1 F0_11_13 ( .D(\din[13][11] ), .G(n73), .Q(\q[13][11] ) );
    LD1 F0_14_2 ( .D(\din[2][14] ), .G(n73), .Q(\q[2][14] ) );
    LD1 F0_9_10 ( .D(\din[10][9] ), .G(n73), .Q(\q[10][9] ) );
    LD1 F0_11_4 ( .D(\din[4][11] ), .G(n73), .Q(\q[4][11] ) );
    LD1 F0_5_13 ( .D(\din[13][5] ), .G(n73), .Q(\q[13][5] ) );
    LD1 F0_3_0 ( .D(\din[0][3] ), .G(n73), .Q(\q[0][3] ) );
    LD1 F0_13_8 ( .D(\din[8][13] ), .G(n73), .Q(\q[8][13] ) );
    LD1 F0_15_2 ( .D(\din[2][15] ), .G(n73), .Q(\q[2][15] ) );
    LD1 F0_10_4 ( .D(\din[4][10] ), .G(n73), .Q(\q[4][10] ) );
    LD1 F0_6_6 ( .D(\din[6][6] ), .G(n73), .Q(\q[6][6] ) );
    LD1 F0_10_12 ( .D(\din[12][10] ), .G(n73), .Q(\q[12][10] ) );
    LD1 F0_7_6 ( .D(\din[6][7] ), .G(n73), .Q(\q[6][7] ) );
    LD1 F0_12_8 ( .D(\din[8][12] ), .G(n73), .Q(\q[8][12] ) );
    LD1 F0_8_11 ( .D(\din[11][8] ), .G(n73), .Q(\q[11][8] ) );
    LD1 F0_4_12 ( .D(\din[12][4] ), .G(n73), .Q(\q[12][4] ) );
    LD1 F0_2_0 ( .D(\din[0][2] ), .G(n73), .Q(\q[0][2] ) );
    LD1 F0_9_4 ( .D(\din[4][9] ), .G(n73), .Q(\q[4][9] ) );
    LD1 F0_1_12 ( .D(\din[12][1] ), .G(n73), .Q(\q[12][1] ) );
    LD1 F0_15_12 ( .D(\din[12][15] ), .G(n73), .Q(\q[12][15] ) );
    LD1 F0_13_1 ( .D(\din[1][13] ), .G(n73), .Q(\q[1][13] ) );
    LD1 F0_4_3 ( .D(\din[3][4] ), .G(n73), .Q(\q[3][4] ) );
    LD1 F0_5_3 ( .D(\din[3][5] ), .G(n73), .Q(\q[3][5] ) );
    LD1 F0_3_9 ( .D(\din[9][3] ), .G(n73), .Q(\q[9][3] ) );
    LD1 F0_1_5 ( .D(\din[5][1] ), .G(n73), .Q(\q[5][1] ) );
    LD1 F0_0_13 ( .D(\din[13][0] ), .G(n73), .Q(\q[13][0] ) );
    LD1 F0_14_13 ( .D(\din[13][14] ), .G(n73), .Q(\q[13][14] ) );
    LD1 F0_12_1 ( .D(\din[1][12] ), .G(n73), .Q(\q[1][12] ) );
    LD1 F0_8_4 ( .D(\din[4][8] ), .G(n73), .Q(\q[4][8] ) );
    LD1 F0_12_11 ( .D(\din[11][12] ), .G(n73), .Q(\q[11][12] ) );
    LD1 F0_8_3 ( .D(\din[3][8] ), .G(n73), .Q(\q[3][8] ) );
    LD1 F0_6_11 ( .D(\din[11][6] ), .G(n73), .Q(\q[11][6] ) );
    LD1 F0_2_9 ( .D(\din[9][2] ), .G(n73), .Q(\q[9][2] ) );
    LD1 F0_14_14 ( .D(\din[14][14] ), .G(n73), .Q(\q[14][14] ) );
    LD1 F0_0_5 ( .D(\din[5][0] ), .G(n73), .Q(\q[5][0] ) );
    LD1 F0_7_8 ( .D(\din[8][7] ), .G(n73), .Q(\q[8][7] ) );
    LD1 F0_5_4 ( .D(\din[4][5] ), .G(n73), .Q(\q[4][5] ) );
    LD1 F0_13_10 ( .D(\din[10][13] ), .G(n73), .Q(\q[10][13] ) );
    LD1 F0_12_6 ( .D(\din[6][12] ), .G(n73), .Q(\q[6][12] ) );
    LD1 F0_4_4 ( .D(\din[4][4] ), .G(n73), .Q(\q[4][4] ) );
    LD1 F0_7_10 ( .D(\din[10][7] ), .G(n73), .Q(\q[10][7] ) );
    LD1 F0_1_2 ( .D(\din[2][1] ), .G(n73), .Q(\q[2][1] ) );
    LD1 F0_0_14 ( .D(\din[14][0] ), .G(n73), .Q(\q[14][0] ) );
    LD1 F0_13_6 ( .D(\din[6][13] ), .G(n73), .Q(\q[6][13] ) );
    LD1 F0_15_15 ( .D(\din[15][15] ), .G(n73), .Q(\q[15][15] ) );
    LD1 F0_6_8 ( .D(\din[8][6] ), .G(n73), .Q(\q[8][6] ) );
    LD1 F0_9_3 ( .D(\din[3][9] ), .G(n73), .Q(\q[3][9] ) );
    LD1 F0_15_5 ( .D(\din[5][15] ), .G(n73), .Q(\q[5][15] ) );
    LD1 F0_10_3 ( .D(\din[3][10] ), .G(n73), .Q(\q[3][10] ) );
    LD1 F0_4_15 ( .D(\din[15][4] ), .G(n73), .Q(\q[15][4] ) );
    LD1 F0_2_10 ( .D(\din[10][2] ), .G(n73), .Q(\q[10][2] ) );
    LD1 F0_10_15 ( .D(\din[15][10] ), .G(n73), .Q(\q[15][10] ) );
    LD1 F0_7_1 ( .D(\din[1][7] ), .G(n73), .Q(\q[1][7] ) );
    LD1 F0_14_5 ( .D(\din[5][14] ), .G(n73), .Q(\q[5][14] ) );
    LD1 F0_11_3 ( .D(\din[3][11] ), .G(n73), .Q(\q[3][11] ) );
    LD1 F0_6_1 ( .D(\din[1][6] ), .G(n73), .Q(\q[1][6] ) );
    LD1 F0_3_11 ( .D(\din[11][3] ), .G(n73), .Q(\q[11][3] ) );
    LD1 F0_2_7 ( .D(\din[7][2] ), .G(n73), .Q(\q[7][2] ) );
    LD1 F0_11_14 ( .D(\din[14][11] ), .G(n73), .Q(\q[14][11] ) );
    LD1 F0_5_14 ( .D(\din[14][5] ), .G(n73), .Q(\q[14][5] ) );
    LD1 F0_15_14 ( .D(\din[14][15] ), .G(n73), .Q(\q[14][15] ) );
    LD1 F0_3_7 ( .D(\din[7][3] ), .G(n73), .Q(\q[7][3] ) );
    LD1 F0_1_15 ( .D(\din[15][1] ), .G(n73), .Q(\q[15][1] ) );
    LD1 F0_9_2 ( .D(\din[2][9] ), .G(n73), .Q(\q[2][9] ) );
    LD1 F0_13_11 ( .D(\din[11][13] ), .G(n73), .Q(\q[11][13] ) );
    LD1 F0_4_5 ( .D(\din[5][4] ), .G(n73), .Q(\q[5][4] ) );
    LD1 F0_1_14 ( .D(\din[14][1] ), .G(n73), .Q(\q[14][1] ) );
    LD1 F0_1_3 ( .D(\din[3][1] ), .G(n73), .Q(\q[3][1] ) );
    LD1 F0_13_7 ( .D(\din[7][13] ), .G(n73), .Q(\q[7][13] ) );
    LD1 F0_7_11 ( .D(\din[11][7] ), .G(n73), .Q(\q[11][7] ) );
    LD1 F0_6_9 ( .D(\din[9][6] ), .G(n73), .Q(\q[9][6] ) );
    LD1 F0_14_15 ( .D(\din[15][14] ), .G(n73), .Q(\q[15][14] ) );
    LD1 F0_12_7 ( .D(\din[7][12] ), .G(n73), .Q(\q[7][12] ) );
    LD1 F0_7_9 ( .D(\din[9][7] ), .G(n73), .Q(\q[9][7] ) );
    LD1 F0_5_5 ( .D(\din[5][5] ), .G(n73), .Q(\q[5][5] ) );
    LD1 F0_12_10 ( .D(\din[10][12] ), .G(n73), .Q(\q[10][12] ) );
    LD1 F0_8_2 ( .D(\din[2][8] ), .G(n73), .Q(\q[2][8] ) );
    LD1 F0_6_10 ( .D(\din[10][6] ), .G(n73), .Q(\q[10][6] ) );
    LD1 F0_11_15 ( .D(\din[15][11] ), .G(n73), .Q(\q[15][11] ) );
    LD1 F0_5_15 ( .D(\din[15][5] ), .G(n73), .Q(\q[15][5] ) );
    LD1 F0_14_4 ( .D(\din[4][14] ), .G(n73), .Q(\q[4][14] ) );
    LD1 F0_11_2 ( .D(\din[2][11] ), .G(n73), .Q(\q[2][11] ) );
    LD1 F0_6_0 ( .D(\din[0][6] ), .G(n73), .Q(\q[0][6] ) );
    LD1 F0_3_10 ( .D(\din[10][3] ), .G(n73), .Q(\q[10][3] ) );
    LD1 F0_3_6 ( .D(\din[6][3] ), .G(n73), .Q(\q[6][3] ) );
    LD1 F0_15_4 ( .D(\din[4][15] ), .G(n73), .Q(\q[4][15] ) );
    LD1 F0_10_2 ( .D(\din[2][10] ), .G(n73), .Q(\q[2][10] ) );
    LD1 F0_4_14 ( .D(\din[14][4] ), .G(n73), .Q(\q[14][4] ) );
    LD1 F0_7_0 ( .D(\din[0][7] ), .G(n73), .Q(\q[0][7] ) );
    LD1 F0_10_14 ( .D(\din[14][10] ), .G(n73), .Q(\q[14][10] ) );
    LD1 F0_15_3 ( .D(\din[3][15] ), .G(n73), .Q(\q[3][15] ) );
    LD1 F0_10_13 ( .D(\din[13][10] ), .G(n73), .Q(\q[13][10] ) );
    LD1 F0_10_5 ( .D(\din[5][10] ), .G(n73), .Q(\q[5][10] ) );
    LD1 F0_8_10 ( .D(\din[10][8] ), .G(n73), .Q(\q[10][8] ) );
    LD1 F0_12_9 ( .D(\din[9][12] ), .G(n73), .Q(\q[9][12] ) );
    LD1 F0_7_7 ( .D(\din[7][7] ), .G(n73), .Q(\q[7][7] ) );
    LD1 F0_2_11 ( .D(\din[11][2] ), .G(n73), .Q(\q[11][2] ) );
    LD1 F0_2_6 ( .D(\din[6][2] ), .G(n73), .Q(\q[6][2] ) );
    LD1 F0_14_3 ( .D(\din[3][14] ), .G(n73), .Q(\q[3][14] ) );
    LD1 F0_9_11 ( .D(\din[11][9] ), .G(n73), .Q(\q[11][9] ) );
    LD1 F0_11_5 ( .D(\din[5][11] ), .G(n73), .Q(\q[5][11] ) );
    LD1 F0_4_13 ( .D(\din[13][4] ), .G(n73), .Q(\q[13][4] ) );
    LD1 F0_13_9 ( .D(\din[9][13] ), .G(n73), .Q(\q[9][13] ) );
    LD1 F0_3_1 ( .D(\din[1][3] ), .G(n73), .Q(\q[1][3] ) );
    LD1 F0_6_7 ( .D(\din[7][6] ), .G(n73), .Q(\q[7][6] ) );
    LD1 F0_11_12 ( .D(\din[12][11] ), .G(n73), .Q(\q[12][11] ) );
    LD1 F0_8_5 ( .D(\din[5][8] ), .G(n73), .Q(\q[5][8] ) );
    LD1 F0_5_12 ( .D(\din[12][5] ), .G(n73), .Q(\q[12][5] ) );
    LD1 F0_5_2 ( .D(\din[2][5] ), .G(n73), .Q(\q[2][5] ) );
    LD1 F0_2_1 ( .D(\din[1][2] ), .G(n73), .Q(\q[1][2] ) );
    LD1 F0_0_15 ( .D(\din[15][0] ), .G(n73), .Q(\q[15][0] ) );
    LD1 F0_14_12 ( .D(\din[12][14] ), .G(n73), .Q(\q[12][14] ) );
    LD1 F0_0_12 ( .D(\din[12][0] ), .G(n73), .Q(\q[12][0] ) );
    LD1 F0_12_0 ( .D(\din[0][12] ), .G(n73), .Q(\q[0][12] ) );
    LD1 F0_2_8 ( .D(\din[8][2] ), .G(n73), .Q(\q[8][2] ) );
    LD1 F0_0_4 ( .D(\din[4][0] ), .G(n73), .Q(\q[4][0] ) );
    LD1 F0_0_3 ( .D(\din[3][0] ), .G(n73), .Q(\q[3][0] ) );
    LD1 F0_13_0 ( .D(\din[0][13] ), .G(n73), .Q(\q[0][13] ) );
    LD1 F0_4_2 ( .D(\din[2][4] ), .G(n73), .Q(\q[2][4] ) );
    LD1 F0_3_8 ( .D(\din[8][3] ), .G(n73), .Q(\q[8][3] ) );
    LD1 F0_9_5 ( .D(\din[5][9] ), .G(n73), .Q(\q[5][9] ) );
    LD1 F0_1_13 ( .D(\din[13][1] ), .G(n73), .Q(\q[13][1] ) );
    LD1 F0_1_4 ( .D(\din[4][1] ), .G(n73), .Q(\q[4][1] ) );
    LD1 F0_15_13 ( .D(\din[13][15] ), .G(n73), .Q(\q[13][15] ) );
    LD1 F0_5_10 ( .D(\din[10][5] ), .G(n73), .Q(\q[10][5] ) );
    LD1 F0_11_10 ( .D(\din[10][11] ), .G(n73), .Q(\q[10][11] ) );
    LD1 F0_6_5 ( .D(\din[5][6] ), .G(n73), .Q(\q[5][6] ) );
    LD1 F0_3_15 ( .D(\din[15][3] ), .G(n73), .Q(\q[15][3] ) );
    LD1 F0_3_3 ( .D(\din[3][3] ), .G(n73), .Q(\q[3][3] ) );
    LD1 F0_11_7 ( .D(\din[7][11] ), .G(n73), .Q(\q[7][11] ) );
    LD1 F0_9_13 ( .D(\din[13][9] ), .G(n73), .Q(\q[13][9] ) );
    LD1 F0_14_1 ( .D(\din[1][14] ), .G(n73), .Q(\q[1][14] ) );
    LD1 F0_4_9 ( .D(\din[9][4] ), .G(n73), .Q(\q[9][4] ) );
    LD1 F0_4_11 ( .D(\din[11][4] ), .G(n73), .Q(\q[11][4] ) );
    LD1 F0_10_11 ( .D(\din[11][10] ), .G(n73), .Q(\q[11][10] ) );
    LD1 F0_7_5 ( .D(\din[5][7] ), .G(n73), .Q(\q[5][7] ) );
    LD1 F0_15_1 ( .D(\din[1][15] ), .G(n73), .Q(\q[1][15] ) );
    LD1 F0_10_7 ( .D(\din[7][10] ), .G(n73), .Q(\q[7][10] ) );
    LD1 F0_5_9 ( .D(\din[9][5] ), .G(n73), .Q(\q[9][5] ) );
    LD1 F0_2_3 ( .D(\din[3][2] ), .G(n73), .Q(\q[3][2] ) );
    LD1 F0_8_12 ( .D(\din[12][8] ), .G(n73), .Q(\q[12][8] ) );
    LD1 F0_2_14 ( .D(\din[14][2] ), .G(n73), .Q(\q[14][2] ) );
    LD1 F0_15_11 ( .D(\din[11][15] ), .G(n73), .Q(\q[11][15] ) );
    LD1 F0_13_2 ( .D(\din[2][13] ), .G(n73), .Q(\q[2][13] ) );
    LD1 F0_9_7 ( .D(\din[7][9] ), .G(n73), .Q(\q[7][9] ) );
    LD1 F0_14_8 ( .D(\din[8][14] ), .G(n73), .Q(\q[8][14] ) );
    LD1 F0_13_14 ( .D(\din[14][13] ), .G(n73), .Q(\q[14][13] ) );
    LD1 F0_4_0 ( .D(\din[0][4] ), .G(n73), .Q(\q[0][4] ) );
    LD1 F0_1_11 ( .D(\din[11][1] ), .G(n73), .Q(\q[11][1] ) );
    LD1 F0_0_2 ( .D(\din[2][0] ), .G(n73), .Q(\q[2][0] ) );
    LD1 F0_7_14 ( .D(\din[14][7] ), .G(n73), .Q(\q[14][7] ) );
    LD1 F0_12_2 ( .D(\din[2][12] ), .G(n73), .Q(\q[2][12] ) );
    LD1 F0_1_6 ( .D(\din[6][1] ), .G(n73), .Q(\q[6][1] ) );
    LD1 F0_14_10 ( .D(\din[10][14] ), .G(n73), .Q(\q[10][14] ) );
    LD1 F0_5_0 ( .D(\din[0][5] ), .G(n73), .Q(\q[0][5] ) );
    LD1 F0_15_8 ( .D(\din[8][15] ), .G(n73), .Q(\q[8][15] ) );
    LD1 F0_12_15 ( .D(\din[15][12] ), .G(n73), .Q(\q[15][12] ) );
    LD1 F0_8_7 ( .D(\din[7][8] ), .G(n73), .Q(\q[7][8] ) );
    LD1 F0_6_15 ( .D(\din[15][6] ), .G(n73), .Q(\q[15][6] ) );
    LD1 F0_12_12 ( .D(\din[12][12] ), .G(n73), .Q(\q[12][12] ) );
    LD1 F0_12_5 ( .D(\din[5][12] ), .G(n73), .Q(\q[5][12] ) );
    LD1 F0_8_0 ( .D(\din[0][8] ), .G(n73), .Q(\q[0][8] ) );
    LD1 F0_6_12 ( .D(\din[12][6] ), .G(n73), .Q(\q[12][6] ) );
    LD1 F0_10_9 ( .D(\din[9][10] ), .G(n73), .Q(\q[9][10] ) );
    LD1 F0_5_7 ( .D(\din[7][5] ), .G(n73), .Q(\q[7][5] ) );
    LD1 F0_0_10 ( .D(\din[10][0] ), .G(n73), .Q(\q[10][0] ) );
    LD1 F0_0_6 ( .D(\din[6][0] ), .G(n73), .Q(\q[6][0] ) );
    LD1 F0_13_5 ( .D(\din[5][13] ), .G(n73), .Q(\q[5][13] ) );
    LD1 F0_11_9 ( .D(\din[9][11] ), .G(n73), .Q(\q[9][11] ) );
    LD1 F0_7_13 ( .D(\din[13][7] ), .G(n73), .Q(\q[13][7] ) );
    LD1 F0_1_1 ( .D(\din[1][1] ), .G(n73), .Q(\q[1][1] ) );
    LD1 F0_13_13 ( .D(\din[13][13] ), .G(n73), .Q(\q[13][13] ) );
    LD1 F0_9_0 ( .D(\din[0][9] ), .G(n73), .Q(\q[0][9] ) );
    LD1 F0_4_7 ( .D(\din[7][4] ), .G(n73), .Q(\q[7][4] ) );
    LD1 F0_8_15 ( .D(\din[15][8] ), .G(n73), .Q(\q[15][8] ) );
    LD1 F0_8_9 ( .D(\din[9][8] ), .G(n73), .Q(\q[9][8] ) );
    LD1 F0_7_2 ( .D(\din[2][7] ), .G(n73), .Q(\q[2][7] ) );
    LD1 F0_2_13 ( .D(\din[13][2] ), .G(n73), .Q(\q[13][2] ) );
    LD1 F0_2_4 ( .D(\din[4][2] ), .G(n73), .Q(\q[4][2] ) );
    LD1 F0_10_0 ( .D(\din[0][10] ), .G(n73), .Q(\q[0][10] ) );
    LD1 F0_15_6 ( .D(\din[6][15] ), .G(n73), .Q(\q[6][15] ) );
    LD1 F0_3_4 ( .D(\din[4][3] ), .G(n73), .Q(\q[4][3] ) );
    LD1 F0_6_2 ( .D(\din[2][6] ), .G(n73), .Q(\q[2][6] ) );
    LD1 F0_14_6 ( .D(\din[6][14] ), .G(n73), .Q(\q[6][14] ) );
    LD1 F0_11_0 ( .D(\din[0][11] ), .G(n73), .Q(\q[0][11] ) );
    LD1 F0_9_14 ( .D(\din[14][9] ), .G(n73), .Q(\q[14][9] ) );
    LD1 F0_3_12 ( .D(\din[12][3] ), .G(n73), .Q(\q[12][3] ) );
    LD1 F0_9_9 ( .D(\din[9][9] ), .G(n73), .Q(\q[9][9] ) );
    LD1 F0_9_1 ( .D(\din[1][9] ), .G(n73), .Q(\q[1][9] ) );
    LD1 F0_13_4 ( .D(\din[4][13] ), .G(n73), .Q(\q[4][13] ) );
    LD1 F0_1_8 ( .D(\din[8][1] ), .G(n73), .Q(\q[8][1] ) );
    LD1 F0_1_0 ( .D(\din[0][1] ), .G(n73), .Q(\q[0][1] ) );
    LD1 F0_0_8 ( .D(\din[8][0] ), .G(n73), .Q(\q[8][0] ) );
    LD1 F0_11_8 ( .D(\din[8][11] ), .G(n73), .Q(\q[8][11] ) );
    LD1 F0_13_12 ( .D(\din[12][13] ), .G(n73), .Q(\q[12][13] ) );
    LD1 F0_7_12 ( .D(\din[12][7] ), .G(n73), .Q(\q[12][7] ) );
    LD1 F0_12_4 ( .D(\din[4][12] ), .G(n73), .Q(\q[4][12] ) );
    LD1 F0_4_6 ( .D(\din[6][4] ), .G(n73), .Q(\q[6][4] ) );
    LD1 F0_5_6 ( .D(\din[6][5] ), .G(n73), .Q(\q[6][5] ) );
    LD1 F0_10_8 ( .D(\din[8][10] ), .G(n73), .Q(\q[8][10] ) );
    LD1 F0_0_1 ( .D(\din[1][0] ), .G(n73), .Q(\q[1][0] ) );
    LD1 F0_12_13 ( .D(\din[13][12] ), .G(n73), .Q(\q[13][12] ) );
    LD1 F0_9_8 ( .D(\din[8][9] ), .G(n73), .Q(\q[8][9] ) );
    LD1 F0_8_1 ( .D(\din[1][8] ), .G(n73), .Q(\q[1][8] ) );
    LD1 F0_6_13 ( .D(\din[13][6] ), .G(n73), .Q(\q[13][6] ) );
    LD1 F0_6_3 ( .D(\din[3][6] ), .G(n73), .Q(\q[3][6] ) );
    LD1 F0_14_7 ( .D(\din[7][14] ), .G(n73), .Q(\q[7][14] ) );
    LD1 F0_11_1 ( .D(\din[1][11] ), .G(n73), .Q(\q[1][11] ) );
    LD1 F0_9_15 ( .D(\din[15][9] ), .G(n73), .Q(\q[15][9] ) );
    LD1 F0_3_13 ( .D(\din[13][3] ), .G(n73), .Q(\q[13][3] ) );
    LD1 F0_3_5 ( .D(\din[5][3] ), .G(n73), .Q(\q[5][3] ) );
    LD1 F0_7_3 ( .D(\din[3][7] ), .G(n73), .Q(\q[3][7] ) );
    LD1 F0_2_5 ( .D(\din[5][2] ), .G(n73), .Q(\q[5][2] ) );
    LD1 F0_1_9 ( .D(\din[9][1] ), .G(n73), .Q(\q[9][1] ) );
    LD1 F0_15_7 ( .D(\din[7][15] ), .G(n73), .Q(\q[7][15] ) );
    LD1 F0_10_1 ( .D(\din[1][10] ), .G(n73), .Q(\q[1][10] ) );
    LD1 F0_8_14 ( .D(\din[14][8] ), .G(n73), .Q(\q[14][8] ) );
    LD1 F0_8_8 ( .D(\din[8][8] ), .G(n73), .Q(\q[8][8] ) );
    LD1 F0_8_13 ( .D(\din[13][8] ), .G(n73), .Q(\q[13][8] ) );
    LD1 F0_4_10 ( .D(\din[10][4] ), .G(n73), .Q(\q[10][4] ) );
    LD1 F0_2_15 ( .D(\din[15][2] ), .G(n73), .Q(\q[15][2] ) );
    LD1 F0_2_12 ( .D(\din[12][2] ), .G(n73), .Q(\q[12][2] ) );
    LD1 F0_10_10 ( .D(\din[10][10] ), .G(n73), .Q(\q[10][10] ) );
    LD1 F0_15_0 ( .D(\din[0][15] ), .G(n73), .Q(\q[0][15] ) );
    LD1 F0_7_4 ( .D(\din[4][7] ), .G(n73), .Q(\q[4][7] ) );
    LD1 F0_5_8 ( .D(\din[8][5] ), .G(n73), .Q(\q[8][5] ) );
    LD1 F0_2_2 ( .D(\din[2][2] ), .G(n73), .Q(\q[2][2] ) );
    LD1 F0_10_6 ( .D(\din[6][10] ), .G(n73), .Q(\q[6][10] ) );
    LD1 F0_6_4 ( .D(\din[4][6] ), .G(n73), .Q(\q[4][6] ) );
    LD1 F0_3_14 ( .D(\din[14][3] ), .G(n73), .Q(\q[14][3] ) );
    LD1 F0_3_2 ( .D(\din[2][3] ), .G(n73), .Q(\q[2][3] ) );
    LD1 F0_0_9 ( .D(\din[9][0] ), .G(n73), .Q(\q[9][0] ) );
    LD1 F0_11_6 ( .D(\din[6][11] ), .G(n73), .Q(\q[6][11] ) );
    LD1 F0_14_0 ( .D(\din[0][14] ), .G(n73), .Q(\q[0][14] ) );
    LD1 F0_9_12 ( .D(\din[12][9] ), .G(n73), .Q(\q[12][9] ) );
    LD1 F0_5_11 ( .D(\din[11][5] ), .G(n73), .Q(\q[11][5] ) );
    LD1 F0_11_11 ( .D(\din[11][11] ), .G(n73), .Q(\q[11][11] ) );
    LD1 F0_12_14 ( .D(\din[14][12] ), .G(n73), .Q(\q[14][12] ) );
    LD1 F0_8_6 ( .D(\din[6][8] ), .G(n73), .Q(\q[6][8] ) );
    LD1 F0_14_11 ( .D(\din[11][14] ), .G(n73), .Q(\q[11][14] ) );
    LD1 F0_12_3 ( .D(\din[3][12] ), .G(n73), .Q(\q[3][12] ) );
    LD1 F0_6_14 ( .D(\din[14][6] ), .G(n73), .Q(\q[14][6] ) );
    LD1 F0_4_8 ( .D(\din[8][4] ), .G(n73), .Q(\q[8][4] ) );
    LD1 F0_15_9 ( .D(\din[9][15] ), .G(n73), .Q(\q[9][15] ) );
    LD1 F0_5_1 ( .D(\din[1][5] ), .G(n73), .Q(\q[1][5] ) );
    LD1 F0_14_9 ( .D(\din[9][14] ), .G(n73), .Q(\q[9][14] ) );
    LD1 F0_13_3 ( .D(\din[3][13] ), .G(n73), .Q(\q[3][13] ) );
    LD1 F0_13_15 ( .D(\din[15][13] ), .G(n73), .Q(\q[15][13] ) );
    LD1 F0_7_15 ( .D(\din[15][7] ), .G(n73), .Q(\q[15][7] ) );
    LD1 F0_4_1 ( .D(\din[1][4] ), .G(n73), .Q(\q[1][4] ) );
    LD1 F0_0_11 ( .D(\din[11][0] ), .G(n73), .Q(\q[11][0] ) );
    LD1 F0_0_7 ( .D(\din[7][0] ), .G(n73), .Q(\q[7][0] ) );
    LD1 F0_0_0 ( .D(\din[0][0] ), .G(n73), .Q(\q[0][0] ) );
    LD1 F0_1_7 ( .D(\din[7][1] ), .G(n73), .Q(\q[7][1] ) );
    LD1 F0_15_10 ( .D(\din[10][15] ), .G(n73), .Q(\q[10][15] ) );
    LD1 F0_9_6 ( .D(\din[6][9] ), .G(n73), .Q(\q[6][9] ) );
    LD1 F0_1_10 ( .D(\din[10][1] ), .G(n73), .Q(\q[10][1] ) );
    NR2 U39 ( .A(n74), .B(wr_n), .Z(\wren[6] ) );
    NR2 U40 ( .A(n75), .B(wr_n), .Z(\wren[1] ) );
    NR2 U41 ( .A(n76), .B(wr_n), .Z(\wren[8] ) );
    NR2 U42 ( .A(n77), .B(wr_n), .Z(\wren[10] ) );
    NR2 U43 ( .A(n78), .B(wr_n), .Z(\wren[0] ) );
    NR2 U44 ( .A(n79), .B(wr_n), .Z(\wren[11] ) );
    NR2 U45 ( .A(n80), .B(wr_n), .Z(\wren[9] ) );
    NR2 U46 ( .A(n81), .B(wr_n), .Z(\wren[7] ) );
    NR2 U47 ( .A(n82), .B(wr_n), .Z(\wren[14] ) );
    NR2 U48 ( .A(n83), .B(wr_n), .Z(\wren[5] ) );
    NR2 U49 ( .A(n84), .B(wr_n), .Z(\wren[2] ) );
    NR2 U50 ( .A(n85), .B(wr_n), .Z(\wren[13] ) );
    NR2 U51 ( .A(n86), .B(wr_n), .Z(\wren[3] ) );
    NR2 U52 ( .A(n87), .B(wr_n), .Z(\wren[12] ) );
    NR2 U53 ( .A(n88), .B(wr_n), .Z(\wren[15] ) );
    NR2 U54 ( .A(n89), .B(wr_n), .Z(\wren[4] ) );
    IV U55 ( .A(clk), .Z(n73) );
    IV U56 ( .A(wr_addr[9]), .Z(n80) );
    IV U57 ( .A(wr_addr[8]), .Z(n76) );
    IV U58 ( .A(wr_addr[7]), .Z(n81) );
    IV U59 ( .A(wr_addr[6]), .Z(n74) );
    IV U60 ( .A(wr_addr[5]), .Z(n83) );
    IV U61 ( .A(wr_addr[4]), .Z(n89) );
    IV U62 ( .A(wr_addr[3]), .Z(n86) );
    IV U63 ( .A(wr_addr[2]), .Z(n84) );
    IV U64 ( .A(wr_addr[1]), .Z(n75) );
    IV U65 ( .A(wr_addr[15]), .Z(n88) );
    IV U66 ( .A(wr_addr[14]), .Z(n82) );
    IV U67 ( .A(wr_addr[13]), .Z(n85) );
    IV U68 ( .A(wr_addr[12]), .Z(n87) );
    IV U69 ( .A(wr_addr[11]), .Z(n79) );
    IV U70 ( .A(wr_addr[10]), .Z(n77) );
    IV U71 ( .A(wr_addr[0]), .Z(n78) );
endmodule


module fifo_DW_ram_r_w_s_lat_32_16_0 ( clk, cs_n, wr_n, rd_addr, wr_addr, 
    data_in, data_out );
output [31:0] data_out;
input  [3:0] rd_addr;
input  [3:0] wr_addr;
input  [31:0] data_in;
input  clk, cs_n, wr_n;
    wire \addr_dec[13] , \addr_dec[15] , \addr_dec[11] , \addr_dec[4] , 
        \addr_dec[0] , \addr_dec[9] , \addr_dec[2] , \addr_dec[6] , 
        \addr_dec[7] , \addr_dec[3] , \addr_dec[1] , \addr_dec[8] , 
        \addr_dec[5] , \addr_dec[10] , \addr_dec[14] , \addr_dec[12] , n90, 
        n91, n92, n94, n95, n96, n97, n98, n99, n100, n101;
    fifo_DW_MEM_R_W_S_LAT_16_16_1 M0_2 ( .clk(clk), .wr_n(wr_n), .rd_addr(
        rd_addr), .wr_addr({\addr_dec[15] , \addr_dec[14] , \addr_dec[13] , 
        \addr_dec[12] , \addr_dec[11] , \addr_dec[10] , \addr_dec[9] , 
        \addr_dec[8] , \addr_dec[7] , \addr_dec[6] , \addr_dec[5] , 
        \addr_dec[4] , \addr_dec[3] , \addr_dec[2] , \addr_dec[1] , 
        \addr_dec[0] }), .data_in(data_in[15:0]), .data_out(data_out[15:0]) );
    fifo_DW_MEM_R_W_S_LAT_16_16_0 M0_1 ( .clk(clk), .wr_n(wr_n), .rd_addr(
        rd_addr), .wr_addr({\addr_dec[15] , \addr_dec[14] , \addr_dec[13] , 
        \addr_dec[12] , \addr_dec[11] , \addr_dec[10] , \addr_dec[9] , 
        \addr_dec[8] , \addr_dec[7] , \addr_dec[6] , \addr_dec[5] , 
        \addr_dec[4] , \addr_dec[3] , \addr_dec[2] , \addr_dec[1] , 
        \addr_dec[0] }), .data_in(data_in[31:16]), .data_out(data_out[31:16])
         );
    NR2 U33 ( .A(n90), .B(n91), .Z(\addr_dec[0] ) );
    NR2 U34 ( .A(n92), .B(n94), .Z(\addr_dec[10] ) );
    NR2 U35 ( .A(n95), .B(n94), .Z(\addr_dec[11] ) );
    NR2 U36 ( .A(n92), .B(n96), .Z(\addr_dec[12] ) );
    NR2 U37 ( .A(n95), .B(n96), .Z(\addr_dec[13] ) );
    NR2 U38 ( .A(n92), .B(n97), .Z(\addr_dec[14] ) );
    NR2 U39 ( .A(n95), .B(n97), .Z(\addr_dec[15] ) );
    NR2 U40 ( .A(n90), .B(n98), .Z(\addr_dec[1] ) );
    NR2 U41 ( .A(n91), .B(n94), .Z(\addr_dec[2] ) );
    NR2 U42 ( .A(n98), .B(n94), .Z(\addr_dec[3] ) );
    NR2 U43 ( .A(n91), .B(n96), .Z(\addr_dec[4] ) );
    NR2 U44 ( .A(n98), .B(n96), .Z(\addr_dec[5] ) );
    NR2 U45 ( .A(n97), .B(n91), .Z(\addr_dec[6] ) );
    NR2 U46 ( .A(n98), .B(n97), .Z(\addr_dec[7] ) );
    NR2 U47 ( .A(n90), .B(n92), .Z(\addr_dec[8] ) );
    NR2 U48 ( .A(n95), .B(n90), .Z(\addr_dec[9] ) );
    ND2 U49 ( .A(wr_addr[3]), .B(wr_addr[0]), .Z(n95) );
    ND2 U50 ( .A(n99), .B(n100), .Z(n90) );
    ND2 U51 ( .A(wr_addr[3]), .B(n101), .Z(n92) );
    IV U52 ( .A(wr_addr[1]), .Z(n99) );
    IV U53 ( .A(wr_addr[2]), .Z(n100) );
    OR2 U54 ( .A(n101), .B(wr_addr[3]), .Z(n98) );
    ND2 U55 ( .A(wr_addr[2]), .B(wr_addr[1]), .Z(n97) );
    ND3 U56 ( .A(n92), .B(n95), .C(n98), .Z(n91) );
    ND2 U57 ( .A(wr_addr[2]), .B(n99), .Z(n96) );
    ND2 U58 ( .A(wr_addr[1]), .B(n100), .Z(n94) );
    IV U59 ( .A(wr_addr[0]), .Z(n101) );
endmodule


module gray2bin_COUNT_WIDTH4_2 ( gray_count, bin_count );
input  [3:0] gray_count;
output [3:0] bin_count;
    wire \gray_count[3] ;
    assign \gray_count[3]  = gray_count[3];
    assign bin_count[3] = \gray_count[3] ;
    EO U10 ( .A(gray_count[0]), .B(bin_count[1]), .Z(bin_count[0]) );
    EO U11 ( .A(\gray_count[3] ), .B(gray_count[2]), .Z(bin_count[2]) );
    EO U12 ( .A(gray_count[1]), .B(bin_count[2]), .Z(bin_count[1]) );
endmodule


module gray2bin_COUNT_WIDTH4_3 ( gray_count, bin_count );
input  [3:0] gray_count;
output [3:0] bin_count;
    wire \gray_count[3] ;
    assign \gray_count[3]  = gray_count[3];
    assign bin_count[3] = \gray_count[3] ;
    EO U10 ( .A(gray_count[0]), .B(bin_count[1]), .Z(bin_count[0]) );
    EO U11 ( .A(\gray_count[3] ), .B(gray_count[2]), .Z(bin_count[2]) );
    EO U12 ( .A(gray_count[1]), .B(bin_count[2]), .Z(bin_count[1]) );
endmodule


module rs_flop_test_1 ( clk, reset_n, s, r, q_out, test_si, test_se );
input  [0:0] s;
output [0:0] q_out;
input  [0:0] r;
input  clk, reset_n, test_si, test_se;
    wire n112, n126, n127;
    FD1S \q_out_reg[0]  ( .D(n112), .CP(clk), .TI(test_si), .TE(test_se), .Q(
        q_out) );
    NR3 U11 ( .A(n126), .B(r), .C(n127), .Z(n112) );
    NR2 U12 ( .A(s), .B(q_out), .Z(n127) );
    IV U13 ( .A(reset_n), .Z(n126) );
endmodule


module gray_counter_WIDTH4_test_2 ( clk, reset, clear, enable, nxt_bin_count, 
    bin_count, gray_count, test_si, test_so, test_se );
output [3:0] nxt_bin_count;
output [3:0] gray_count;
output [3:0] bin_count;
input  clk, reset, clear, enable, test_si, test_se;
output test_so;
    wire test_so_wire, n204, n208, n211, n215, n219, n223, n227, n231, n235, 
        n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
        n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
        n260, n261, n262, n263, n264;
    assign gray_count[3] = test_so_wire;
    assign test_so = test_so_wire;
    FD1S \bin_count_reg[0]  ( .D(n211), .CP(clk), .TI(test_si), .TE(test_se), 
        .Q(bin_count[0]), .QN(n264) );
    FD1S \bin_count_reg[1]  ( .D(n215), .CP(clk), .TI(bin_count[0]), .TE(
        test_se), .Q(bin_count[1]), .QN(n263) );
    FD1S \bin_count_reg[2]  ( .D(n219), .CP(clk), .TI(bin_count[1]), .TE(
        test_se), .Q(bin_count[2]), .QN(n262) );
    FD1S \bin_count_reg[3]  ( .D(n223), .CP(clk), .TI(bin_count[2]), .TE(
        test_se), .Q(bin_count[3]), .QN(n261) );
    FD1S \prsnt_state_reg[3]  ( .D(n208), .CP(clk), .TI(gray_count[2]), .TE(
        test_se), .Q(test_so_wire), .QN(n235) );
    FD1S \prsnt_state_reg[2]  ( .D(n204), .CP(clk), .TI(gray_count[1]), .TE(
        test_se), .Q(gray_count[2]), .QN(n236) );
    FD1S \prsnt_state_reg[1]  ( .D(n231), .CP(clk), .TI(gray_count[0]), .TE(
        test_se), .Q(gray_count[1]), .QN(n237) );
    FD1S \prsnt_state_reg[0]  ( .D(n227), .CP(clk), .TI(bin_count[3]), .TE(
        test_se), .Q(gray_count[0]), .QN(n238) );
    AO4 U77 ( .A(n236), .B(n239), .C(n240), .D(n241), .Z(n204) );
    AO4 U78 ( .A(n241), .B(n242), .C(n235), .D(n239), .Z(n208) );
    AO4 U79 ( .A(n241), .B(n243), .C(n239), .D(n264), .Z(n211) );
    AO4 U80 ( .A(n244), .B(n241), .C(n239), .D(n263), .Z(n215) );
    AO4 U81 ( .A(n245), .B(n241), .C(n239), .D(n262), .Z(n219) );
    AO4 U82 ( .A(n241), .B(n242), .C(n239), .D(n261), .Z(n223) );
    AO4 U83 ( .A(n238), .B(n239), .C(n246), .D(n241), .Z(n227) );
    AO4 U84 ( .A(n237), .B(n239), .C(n247), .D(n241), .Z(n231) );
    AO2 U85 ( .A(nxt_bin_count[1]), .B(n248), .C(nxt_bin_count[2]), .D(n249), 
        .Z(n247) );
    EO1 U86 ( .A(nxt_bin_count[0]), .B(n249), .C(n244), .D(n250), .Z(n246) );
    AO2 U87 ( .A(nxt_bin_count[3]), .B(n248), .C(n251), .D(nxt_bin_count[2]), 
        .Z(n240) );
    AO4 U88 ( .A(n235), .B(n236), .C(test_so_wire), .D(gray_count[2]), .Z(n252
        ) );
    AO4 U89 ( .A(n254), .B(n237), .C(n252), .D(gray_count[1]), .Z(n253) );
    AO4 U90 ( .A(n238), .B(n255), .C(gray_count[0]), .D(n253), .Z(n250) );
    EO1 U91 ( .A(test_so_wire), .B(n256), .C(test_so_wire), .D(n256), .Z(n251)
         );
    EO1 U92 ( .A(n252), .B(n257), .C(n252), .D(n257), .Z(n248) );
    AO2 U93 ( .A(n255), .B(n258), .C(n253), .D(n259), .Z(n249) );
    IV U94 ( .A(enable), .Z(n260) );
    NR2 U95 ( .A(n260), .B(n250), .Z(n258) );
    NR2 U96 ( .A(n259), .B(n255), .Z(n257) );
    NR2 U97 ( .A(n249), .B(clear), .Z(nxt_bin_count[1]) );
    NR2 U98 ( .A(n248), .B(clear), .Z(nxt_bin_count[2]) );
    ND2 U99 ( .A(reset), .B(enable), .Z(n241) );
    ND2 U100 ( .A(reset), .B(n260), .Z(n239) );
    AO1 U101 ( .A(n260), .B(n250), .C(n258), .D(clear), .Z(nxt_bin_count[0])
         );
    NR2 U102 ( .A(n251), .B(clear), .Z(nxt_bin_count[3]) );
    IV U103 ( .A(nxt_bin_count[2]), .Z(n245) );
    IV U104 ( .A(nxt_bin_count[1]), .Z(n244) );
    IV U105 ( .A(nxt_bin_count[3]), .Z(n242) );
    ND2 U106 ( .A(n257), .B(n254), .Z(n256) );
    IV U107 ( .A(nxt_bin_count[0]), .Z(n243) );
    IV U108 ( .A(n252), .Z(n254) );
    IV U109 ( .A(n253), .Z(n255) );
    IV U110 ( .A(n258), .Z(n259) );
endmodule


module push_ctrl_DEPTH16_counter_width4_almost_full_level8_test_1 ( push_clk, 
    reset_n, pop_count, push, push_full, almost_full, bin_count, push_count, 
    test_si, test_se );
input  [3:0] pop_count;
output [3:0] bin_count;
output [3:0] push_count;
input  push_clk, reset_n, push, test_si, test_se;
output push_full, almost_full;
    wire \pop_count_svd56[0] , \nxt_push_count[1] , \sync_pop_count[0] , 
        \sync_pop_count49[1] , count_enable, \sync_pop_count49[3] , 
        \sync_pop_count[2] , \nxt_push_count[3] , \pop_count_svd56[2] , 
        \sync_pop_countb[1] , \pop_count_svd[3] , counter_clear, 
        \pop_count_svdb[0] , \sync_pop_countb[3] , \pop_count_svd[1] , 
        \sync_pop_countb[2] , \pop_count_svd[0] , \pop_count_svd[2] , 
        \sync_pop_countb[0] , \sync_pop_count[3] , \nxt_push_count[2] , 
        make_full, internal_pop, \pop_count_svd56[3] , \sync_pop_count49[2] , 
        \sync_pop_count49[0] , \pop_count_svd56[1] , \nxt_push_count[0] , 
        \sync_pop_count[1] , n157, n158, n159, n160, n202, n265, n266, n267, 
        n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279;
    wire SYNOPSYS_UNCONNECTED_1 , SYNOPSYS_UNCONNECTED_2 , 
	SYNOPSYS_UNCONNECTED_3 ;
    gray2bin_COUNT_WIDTH4_3 synch1 ( .gray_count({\sync_pop_count[3] , 
        \sync_pop_count[2] , \sync_pop_count[1] , \sync_pop_count[0] }), 
        .bin_count({\sync_pop_countb[3] , \sync_pop_countb[2] , 
        \sync_pop_countb[1] , \sync_pop_countb[0] }) );
    gray2bin_COUNT_WIDTH4_2 synch2 ( .gray_count({\pop_count_svd[3] , 
        \pop_count_svd[2] , \pop_count_svd[1] , \pop_count_svd[0] }), 
        .bin_count({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, \pop_count_svdb[0] }) );
    rs_flop_test_1 full_flag ( .clk(push_clk), .reset_n(reset_n), .s(make_full
        ), .r(internal_pop), .q_out(push_full), .test_si(\sync_pop_count[3] ), 
        .test_se(test_se) );
    gray_counter_WIDTH4_test_2 push_counter ( .clk(push_clk), .reset(reset_n), 
        .clear(counter_clear), .enable(count_enable), .nxt_bin_count({
        \nxt_push_count[3] , \nxt_push_count[2] , \nxt_push_count[1] , 
        \nxt_push_count[0] }), .bin_count(bin_count), .gray_count(push_count), 
        .test_si(\pop_count_svd[3] ), .test_so(n202), .test_se(test_se) );
    FD1S \pop_count_svd_reg[0]  ( .D(\pop_count_svd56[0] ), .CP(push_clk), 
        .TI(test_si), .TE(test_se), .Q(\pop_count_svd[0] ) );
    FD1S \pop_count_svd_reg[1]  ( .D(\pop_count_svd56[1] ), .CP(push_clk), 
        .TI(\pop_count_svd[0] ), .TE(test_se), .Q(\pop_count_svd[1] ) );
    FD1S \pop_count_svd_reg[2]  ( .D(\pop_count_svd56[2] ), .CP(push_clk), 
        .TI(\pop_count_svd[1] ), .TE(test_se), .Q(\pop_count_svd[2] ) );
    FD1S \pop_count_svd_reg[3]  ( .D(\pop_count_svd56[3] ), .CP(push_clk), 
        .TI(\pop_count_svd[2] ), .TE(test_se), .Q(\pop_count_svd[3] ) );
    FD1S \sync_pop_count_reg[0]  ( .D(\sync_pop_count49[0] ), .CP(push_clk), 
        .TI(n202), .TE(test_se), .Q(\sync_pop_count[0] ), .QN(n160) );
    FD1S \sync_pop_count_reg[1]  ( .D(\sync_pop_count49[1] ), .CP(push_clk), 
        .TI(\sync_pop_count[0] ), .TE(test_se), .Q(\sync_pop_count[1] ), .QN(
        n159) );
    FD1S \sync_pop_count_reg[2]  ( .D(\sync_pop_count49[2] ), .CP(push_clk), 
        .TI(\sync_pop_count[1] ), .TE(test_se), .Q(\sync_pop_count[2] ), .QN(
        n158) );
    FD1S \sync_pop_count_reg[3]  ( .D(\sync_pop_count49[3] ), .CP(push_clk), 
        .TI(\sync_pop_count[2] ), .TE(test_se), .Q(\sync_pop_count[3] ), .QN(
        n157) );
    AN2 U43 ( .A(reset_n), .B(pop_count[3]), .Z(\sync_pop_count49[3] ) );
    AN2 U44 ( .A(pop_count[2]), .B(reset_n), .Z(\sync_pop_count49[2] ) );
    AN2 U45 ( .A(pop_count[1]), .B(reset_n), .Z(\sync_pop_count49[1] ) );
    AN2 U46 ( .A(pop_count[0]), .B(reset_n), .Z(\sync_pop_count49[0] ) );
    NR2 U47 ( .A(n265), .B(n157), .Z(\pop_count_svd56[3] ) );
    NR2 U48 ( .A(n265), .B(n158), .Z(\pop_count_svd56[2] ) );
    NR2 U49 ( .A(n265), .B(n159), .Z(\pop_count_svd56[1] ) );
    NR2 U50 ( .A(n265), .B(n160), .Z(\pop_count_svd56[0] ) );
    NR4 U51 ( .A(n266), .B(n267), .C(n268), .D(n269), .Z(make_full) );
    AN4 U52 ( .A(bin_count[3]), .B(bin_count[1]), .C(bin_count[0]), .D(
        bin_count[2]), .Z(counter_clear) );
    AN2 U53 ( .A(n270), .B(push), .Z(count_enable) );
    ND2 U54 ( .A(n271), .B(n270), .Z(almost_full) );
    EO1 U55 ( .A(\sync_pop_countb[0] ), .B(n273), .C(n274), .D(bin_count[1]), 
        .Z(n272) );
    AO6 U56 ( .A(bin_count[1]), .B(n274), .C(n272), .Z(n275) );
    AO5 U57 ( .A(n275), .B(n277), .C(\sync_pop_countb[2] ), .Z(n276) );
    IV U58 ( .A(reset_n), .Z(n265) );
    IV U59 ( .A(\sync_pop_countb[1] ), .Z(n274) );
    IV U60 ( .A(bin_count[2]), .Z(n277) );
    EO U61 ( .A(\nxt_push_count[3] ), .B(\sync_pop_countb[3] ), .Z(n266) );
    EO1 U62 ( .A(\nxt_push_count[1] ), .B(\sync_pop_countb[1] ), .C(
        \nxt_push_count[1] ), .D(\sync_pop_countb[1] ), .Z(n268) );
    EO U63 ( .A(\sync_pop_countb[2] ), .B(\nxt_push_count[2] ), .Z(n269) );
    EO U64 ( .A(\sync_pop_countb[0] ), .B(\pop_count_svdb[0] ), .Z(
        internal_pop) );
    EO U65 ( .A(n276), .B(n278), .Z(n271) );
    ND2 U66 ( .A(n279), .B(push), .Z(n267) );
    EO U67 ( .A(bin_count[3]), .B(\sync_pop_countb[3] ), .Z(n278) );
    IV U68 ( .A(push_full), .Z(n270) );
    EN U69 ( .A(\nxt_push_count[0] ), .B(\sync_pop_countb[0] ), .Z(n279) );
    IV U70 ( .A(bin_count[0]), .Z(n273) );
endmodule


module gray2bin_COUNT_WIDTH4_0 ( gray_count, bin_count );
input  [3:0] gray_count;
output [3:0] bin_count;
    wire \gray_count[3] ;
    assign \gray_count[3]  = gray_count[3];
    assign bin_count[3] = \gray_count[3] ;
    EO U10 ( .A(gray_count[0]), .B(bin_count[1]), .Z(bin_count[0]) );
    EO U11 ( .A(\gray_count[3] ), .B(gray_count[2]), .Z(bin_count[2]) );
    EO U12 ( .A(gray_count[1]), .B(bin_count[2]), .Z(bin_count[1]) );
endmodule


module gray2bin_COUNT_WIDTH4_1 ( gray_count, bin_count );
input  [3:0] gray_count;
output [3:0] bin_count;
    wire \gray_count[3] ;
    assign \gray_count[3]  = gray_count[3];
    assign bin_count[3] = \gray_count[3] ;
    EO U10 ( .A(gray_count[0]), .B(bin_count[1]), .Z(bin_count[0]) );
    EO U11 ( .A(\gray_count[3] ), .B(gray_count[2]), .Z(bin_count[2]) );
    EO U12 ( .A(gray_count[1]), .B(bin_count[2]), .Z(bin_count[1]) );
endmodule


module rs_flop_width1_reset_value1_test_1 ( clk, reset_n, s, r, q_out, test_si, 
    test_se );
input  [0:0] s;
output [0:0] q_out;
input  [0:0] r;
input  clk, reset_n, test_si, test_se;
    wire n91, n93;
    FD1S \q_out_reg[0]  ( .D(n91), .CP(clk), .TI(test_si), .TE(test_se), .Q(
        q_out) );
    AO7 U16 ( .A(r), .B(n93), .C(reset_n), .Z(n91) );
    NR2 U17 ( .A(s), .B(q_out), .Z(n93) );
endmodule


module gray_counter_WIDTH4_test_1 ( clk, reset, clear, enable, nxt_bin_count, 
    bin_count, gray_count, test_si, test_so, test_se );
output [3:0] nxt_bin_count;
output [3:0] gray_count;
output [3:0] bin_count;
input  clk, reset, clear, enable, test_si, test_se;
output test_so;
    wire test_so_wire, n137, n141, n145, n149, n153, n157, n193, n197, n201, 
        n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
        n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, 
        n226, n227, n228, n229, n230;
    assign gray_count[3] = test_so_wire;
    assign test_so = test_so_wire;
    FD1S \bin_count_reg[0]  ( .D(n137), .CP(clk), .TI(test_si), .TE(test_se), 
        .Q(bin_count[0]), .QN(n230) );
    FD1S \bin_count_reg[1]  ( .D(n141), .CP(clk), .TI(bin_count[0]), .TE(
        test_se), .Q(bin_count[1]), .QN(n229) );
    FD1S \bin_count_reg[2]  ( .D(n145), .CP(clk), .TI(bin_count[1]), .TE(
        test_se), .Q(bin_count[2]), .QN(n228) );
    FD1S \bin_count_reg[3]  ( .D(n149), .CP(clk), .TI(bin_count[2]), .TE(
        test_se), .Q(bin_count[3]), .QN(n227) );
    FD1S \prsnt_state_reg[3]  ( .D(n197), .CP(clk), .TI(gray_count[2]), .TE(
        test_se), .Q(test_so_wire), .QN(n201) );
    FD1S \prsnt_state_reg[2]  ( .D(n193), .CP(clk), .TI(gray_count[1]), .TE(
        test_se), .Q(gray_count[2]), .QN(n202) );
    FD1S \prsnt_state_reg[1]  ( .D(n157), .CP(clk), .TI(gray_count[0]), .TE(
        test_se), .Q(gray_count[1]), .QN(n203) );
    FD1S \prsnt_state_reg[0]  ( .D(n153), .CP(clk), .TI(bin_count[3]), .TE(
        test_se), .Q(gray_count[0]), .QN(n204) );
    AO4 U85 ( .A(n205), .B(n206), .C(n207), .D(n230), .Z(n137) );
    AO4 U86 ( .A(n205), .B(n208), .C(n207), .D(n229), .Z(n141) );
    AO4 U87 ( .A(n205), .B(n209), .C(n207), .D(n228), .Z(n145) );
    AO4 U88 ( .A(n205), .B(n210), .C(n207), .D(n227), .Z(n149) );
    AO4 U89 ( .A(n204), .B(n207), .C(n211), .D(n205), .Z(n153) );
    AO4 U90 ( .A(n203), .B(n207), .C(n212), .D(n205), .Z(n157) );
    AO4 U91 ( .A(n202), .B(n207), .C(n213), .D(n205), .Z(n193) );
    AO4 U92 ( .A(n205), .B(n210), .C(n201), .D(n207), .Z(n197) );
    AO2 U93 ( .A(n214), .B(nxt_bin_count[3]), .C(nxt_bin_count[2]), .D(n215), 
        .Z(n213) );
    AO2 U94 ( .A(nxt_bin_count[1]), .B(n214), .C(n216), .D(nxt_bin_count[2]), 
        .Z(n212) );
    EO1 U95 ( .A(nxt_bin_count[0]), .B(n216), .C(n208), .D(n217), .Z(n211) );
    AO4 U96 ( .A(n201), .B(n202), .C(test_so_wire), .D(gray_count[2]), .Z(n218
        ) );
    AO4 U97 ( .A(n220), .B(n203), .C(n218), .D(gray_count[1]), .Z(n219) );
    AO4 U98 ( .A(n204), .B(n221), .C(gray_count[0]), .D(n219), .Z(n217) );
    EO1 U99 ( .A(test_so_wire), .B(n222), .C(test_so_wire), .D(n222), .Z(n215)
         );
    EO1 U100 ( .A(n218), .B(n223), .C(n218), .D(n223), .Z(n214) );
    AO2 U101 ( .A(n221), .B(n224), .C(n219), .D(n225), .Z(n216) );
    IV U102 ( .A(enable), .Z(n226) );
    NR2 U103 ( .A(n226), .B(n217), .Z(n224) );
    NR2 U104 ( .A(n225), .B(n221), .Z(n223) );
    ND2 U105 ( .A(reset), .B(n226), .Z(n207) );
    ND2 U106 ( .A(reset), .B(enable), .Z(n205) );
    NR2 U107 ( .A(n215), .B(clear), .Z(nxt_bin_count[3]) );
    NR2 U108 ( .A(n214), .B(clear), .Z(nxt_bin_count[2]) );
    NR2 U109 ( .A(n216), .B(clear), .Z(nxt_bin_count[1]) );
    AO1 U110 ( .A(n226), .B(n217), .C(n224), .D(clear), .Z(nxt_bin_count[0])
         );
    IV U111 ( .A(nxt_bin_count[2]), .Z(n209) );
    IV U112 ( .A(nxt_bin_count[1]), .Z(n208) );
    IV U113 ( .A(nxt_bin_count[3]), .Z(n210) );
    ND2 U114 ( .A(n223), .B(n220), .Z(n222) );
    IV U115 ( .A(nxt_bin_count[0]), .Z(n206) );
    IV U116 ( .A(n218), .Z(n220) );
    IV U117 ( .A(n219), .Z(n221) );
    IV U118 ( .A(n224), .Z(n225) );
endmodule


module pop_ctrl_DEPTH16_counter_width4_almost_empty_level8_test_1 ( pop_clk, 
    reset_n, push_count, pop, pop_empty, almost_empty, bin_count, pop_count, 
    test_si, test_se );
input  [3:0] push_count;
output [3:0] bin_count;
output [3:0] pop_count;
input  pop_clk, reset_n, pop, test_si, test_se;
output pop_empty, almost_empty;
    wire \push_count_svd56[2] , \sync_push_count49[0] , \sync_push_count[0] , 
        count_enable, \sync_push_count[2] , \sync_push_count49[2] , 
        \push_count_svd56[0] , \nxt_pop_count[0] , \push_count_svd[0] , 
        \sync_push_countb[2] , counter_clear, \sync_push_countb[0] , 
        \push_count_svd[2] , \nxt_pop_count[2] , \push_count_svd[3] , 
        \nxt_pop_count[3] , \sync_push_countb[1] , \sync_push_countb[3] , 
        internal_push, \nxt_pop_count[1] , \push_count_svd[1] , 
        \sync_push_count49[3] , \push_count_svd56[1] , \sync_push_count[3] , 
        \sync_push_count[1] , \push_count_svdb[0] , make_empty, 
        \push_count_svd56[3] , \sync_push_count49[1] , n104, n105, n106, n107, 
        n109, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
        n122, n123, n124, n125;
    wire SYNOPSYS_UNCONNECTED_1 , SYNOPSYS_UNCONNECTED_2 , 
	SYNOPSYS_UNCONNECTED_3 ;
    gray2bin_COUNT_WIDTH4_1 synch1 ( .gray_count({\sync_push_count[3] , 
        \sync_push_count[2] , \sync_push_count[1] , \sync_push_count[0] }), 
        .bin_count({\sync_push_countb[3] , \sync_push_countb[2] , 
        \sync_push_countb[1] , \sync_push_countb[0] }) );
    gray2bin_COUNT_WIDTH4_0 synch2 ( .gray_count({\push_count_svd[3] , 
        \push_count_svd[2] , \push_count_svd[1] , \push_count_svd[0] }), 
        .bin_count({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, \push_count_svdb[0] }) );
    rs_flop_width1_reset_value1_test_1 empty_flag ( .clk(pop_clk), .reset_n(
        reset_n), .s(make_empty), .r(internal_push), .q_out(pop_empty), 
        .test_si(\sync_push_count[3] ), .test_se(test_se) );
    gray_counter_WIDTH4_test_1 push_counter ( .clk(pop_clk), .reset(reset_n), 
        .clear(counter_clear), .enable(count_enable), .nxt_bin_count({
        \nxt_pop_count[3] , \nxt_pop_count[2] , \nxt_pop_count[1] , 
        \nxt_pop_count[0] }), .bin_count(bin_count), .gray_count(pop_count), 
        .test_si(\push_count_svd[3] ), .test_so(n109), .test_se(test_se) );
    FD1S \push_count_svd_reg[0]  ( .D(\push_count_svd56[0] ), .CP(pop_clk), 
        .TI(test_si), .TE(test_se), .Q(\push_count_svd[0] ) );
    FD1S \push_count_svd_reg[1]  ( .D(\push_count_svd56[1] ), .CP(pop_clk), 
        .TI(\push_count_svd[0] ), .TE(test_se), .Q(\push_count_svd[1] ) );
    FD1S \push_count_svd_reg[2]  ( .D(\push_count_svd56[2] ), .CP(pop_clk), 
        .TI(\push_count_svd[1] ), .TE(test_se), .Q(\push_count_svd[2] ) );
    FD1S \push_count_svd_reg[3]  ( .D(\push_count_svd56[3] ), .CP(pop_clk), 
        .TI(\push_count_svd[2] ), .TE(test_se), .Q(\push_count_svd[3] ) );
    FD1S \sync_push_count_reg[0]  ( .D(\sync_push_count49[0] ), .CP(pop_clk), 
        .TI(n109), .TE(test_se), .Q(\sync_push_count[0] ), .QN(n107) );
    FD1S \sync_push_count_reg[1]  ( .D(\sync_push_count49[1] ), .CP(pop_clk), 
        .TI(\sync_push_count[0] ), .TE(test_se), .Q(\sync_push_count[1] ), 
        .QN(n106) );
    FD1S \sync_push_count_reg[2]  ( .D(\sync_push_count49[2] ), .CP(pop_clk), 
        .TI(\sync_push_count[1] ), .TE(test_se), .Q(\sync_push_count[2] ), 
        .QN(n105) );
    FD1S \sync_push_count_reg[3]  ( .D(\sync_push_count49[3] ), .CP(pop_clk), 
        .TI(\sync_push_count[2] ), .TE(test_se), .Q(\sync_push_count[3] ), 
        .QN(n104) );
    AN2 U43 ( .A(reset_n), .B(push_count[3]), .Z(\sync_push_count49[3] ) );
    AN2 U44 ( .A(push_count[2]), .B(reset_n), .Z(\sync_push_count49[2] ) );
    AN2 U45 ( .A(push_count[1]), .B(reset_n), .Z(\sync_push_count49[1] ) );
    AN2 U46 ( .A(push_count[0]), .B(reset_n), .Z(\sync_push_count49[0] ) );
    NR2 U47 ( .A(n111), .B(n104), .Z(\push_count_svd56[3] ) );
    NR2 U48 ( .A(n111), .B(n105), .Z(\push_count_svd56[2] ) );
    NR2 U49 ( .A(n111), .B(n106), .Z(\push_count_svd56[1] ) );
    NR2 U50 ( .A(n111), .B(n107), .Z(\push_count_svd56[0] ) );
    NR4 U51 ( .A(n112), .B(n113), .C(n114), .D(n115), .Z(make_empty) );
    AN4 U52 ( .A(bin_count[3]), .B(bin_count[1]), .C(bin_count[0]), .D(
        bin_count[2]), .Z(counter_clear) );
    AN2 U53 ( .A(n116), .B(pop), .Z(count_enable) );
    ND2 U54 ( .A(n117), .B(n116), .Z(almost_empty) );
    EO1 U55 ( .A(\sync_push_countb[0] ), .B(n119), .C(n120), .D(bin_count[1]), 
        .Z(n118) );
    AO6 U56 ( .A(bin_count[1]), .B(n120), .C(n118), .Z(n121) );
    AO5 U57 ( .A(n121), .B(n123), .C(\sync_push_countb[2] ), .Z(n122) );
    IV U58 ( .A(reset_n), .Z(n111) );
    IV U59 ( .A(\sync_push_countb[1] ), .Z(n120) );
    IV U60 ( .A(bin_count[2]), .Z(n123) );
    EO U61 ( .A(\nxt_pop_count[3] ), .B(\sync_push_countb[3] ), .Z(n112) );
    EO1 U62 ( .A(\nxt_pop_count[1] ), .B(\sync_push_countb[1] ), .C(
        \nxt_pop_count[1] ), .D(\sync_push_countb[1] ), .Z(n114) );
    EO U63 ( .A(\sync_push_countb[2] ), .B(\nxt_pop_count[2] ), .Z(n115) );
    EO U64 ( .A(\sync_push_countb[0] ), .B(\push_count_svdb[0] ), .Z(
        internal_push) );
    EO U65 ( .A(n122), .B(n124), .Z(n117) );
    ND2 U66 ( .A(n125), .B(pop), .Z(n113) );
    EO U67 ( .A(bin_count[3]), .B(\sync_push_countb[3] ), .Z(n124) );
    IV U68 ( .A(pop_empty), .Z(n116) );
    EN U69 ( .A(\nxt_pop_count[0] ), .B(\sync_push_countb[0] ), .Z(n125) );
    IV U70 ( .A(bin_count[0]), .Z(n119) );
endmodule


module fifo ( push_clk, pop_clk, reset_n, push, pop, data_in, data_out, 
    pop_empty, push_full, almost_empty, almost_full, test_si1, test_si2, 
    test_se );
input  [31:0] data_in;
output [31:0] data_out;
input  push_clk, pop_clk, reset_n, push, pop, test_si1, test_si2, test_se;
output pop_empty, push_full, almost_empty, almost_full;
    wire \dataout[6] , \push_count[2] , \dataout[2] , \rd_address[3] , 
        \dataout[9] , \rd_address[1] , \dataout[0] , \push_count[0] , 
        \dataout[4] , \wr_address[0] , \dataout[25] , \dataout[16] , 
        \pop_count[2] , \dataout[21] , \dataout[12] , \dataout[31] , 
        \dataout[28] , \dataout[23] , \dataout[19] , \dataout[10] , 
        \pop_count[0] , \pop_count[1] , \wr_address[2] , \dataout[27] , 
        \dataout[14] , \wr_address[3] , \dataout[26] , \dataout[15] , 
        \dataout[22] , \dataout[18] , \dataout[11] , \dataout[20] , 
        \dataout[13] , \dataout[30] , \dataout[29] , \wr_address[1] , 
        \dataout[24] , \dataout[17] , \pop_count[3] , \push_count[1] , 
        \dataout[5] , \rd_address[0] , \dataout[8] , \dataout[1] , 
        push_clk_inv,
        \dataout[3] , \rd_address[2] , n57, \dataout[7] , \push_count[3] , 
        n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
        n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
        n304, n305, n306, n307, n308, n309, n310, n311;
    fifo_DW_ram_r_w_s_lat_32_16_0 memory ( .clk(push_clk), .cs_n(1'b0), .wr_n(
        n57), .rd_addr({\rd_address[3] , \rd_address[2] , \rd_address[1] , 
        \rd_address[0] }), .wr_addr({\wr_address[3] , \wr_address[2] , 
        \wr_address[1] , \wr_address[0] }), .data_in(data_in), .data_out({
        \dataout[31] , \dataout[30] , \dataout[29] , \dataout[28] , 
        \dataout[27] , \dataout[26] , \dataout[25] , \dataout[24] , 
        \dataout[23] , \dataout[22] , \dataout[21] , \dataout[20] , 
        \dataout[19] , \dataout[18] , \dataout[17] , \dataout[16] , 
        \dataout[15] , \dataout[14] , \dataout[13] , \dataout[12] , 
        \dataout[11] , \dataout[10] , \dataout[9] , \dataout[8] , \dataout[7] , 
        \dataout[6] , \dataout[5] , \dataout[4] , \dataout[3] , \dataout[2] , 
        \dataout[1] , \dataout[0] }) );
    push_ctrl_DEPTH16_counter_width4_almost_full_level8_test_1 push_logic ( 
        .push_clk(push_clk), .reset_n(reset_n), .pop_count({\pop_count[3] , 
        \pop_count[2] , \pop_count[1] , \pop_count[0] }), .push(push), 
        .push_full(push_full), .almost_full(almost_full), .bin_count({
        \wr_address[3] , \wr_address[2] , \wr_address[1] , \wr_address[0] }), 
        .push_count({\push_count[3] , \push_count[2] , \push_count[1] , 
        \push_count[0] }), .test_si(test_si1), .test_se(test_se) );
    pop_ctrl_DEPTH16_counter_width4_almost_empty_level8_test_1 pop_logic ( 
        .pop_clk(pop_clk), .reset_n(reset_n), .push_count({\push_count[3] , 
        \push_count[2] , \push_count[1] , \push_count[0] }), .pop(pop), 
        .pop_empty(pop_empty), .almost_empty(almost_empty), .bin_count({
        \rd_address[3] , \rd_address[2] , \rd_address[1] , \rd_address[0] }), 
        .pop_count({\pop_count[3] , \pop_count[2] , \pop_count[1] , 
        \pop_count[0] }), .test_si(test_si2), .test_se(test_se) );
    IV U81 ( .A(push), .Z(n57) );
    //IV U181 ( .A(push_clk), .Z(push_clk_inv) );
    NR2 U82 ( .A(n280), .B(pop_empty), .Z(data_out[31]) );
    NR2 U83 ( .A(n281), .B(pop_empty), .Z(data_out[30]) );
    NR2 U84 ( .A(n282), .B(pop_empty), .Z(data_out[29]) );
    NR2 U85 ( .A(n283), .B(pop_empty), .Z(data_out[28]) );
    NR2 U86 ( .A(n284), .B(pop_empty), .Z(data_out[27]) );
    NR2 U87 ( .A(n285), .B(pop_empty), .Z(data_out[26]) );
    NR2 U88 ( .A(n286), .B(pop_empty), .Z(data_out[25]) );
    NR2 U89 ( .A(n287), .B(pop_empty), .Z(data_out[24]) );
    NR2 U90 ( .A(n288), .B(pop_empty), .Z(data_out[23]) );
    NR2 U91 ( .A(n289), .B(pop_empty), .Z(data_out[22]) );
    NR2 U92 ( .A(n290), .B(pop_empty), .Z(data_out[21]) );
    NR2 U93 ( .A(n291), .B(pop_empty), .Z(data_out[20]) );
    NR2 U94 ( .A(n292), .B(pop_empty), .Z(data_out[19]) );
    NR2 U95 ( .A(n293), .B(pop_empty), .Z(data_out[18]) );
    NR2 U96 ( .A(n294), .B(pop_empty), .Z(data_out[17]) );
    NR2 U97 ( .A(n295), .B(pop_empty), .Z(data_out[16]) );
    NR2 U98 ( .A(n296), .B(pop_empty), .Z(data_out[15]) );
    NR2 U99 ( .A(n297), .B(pop_empty), .Z(data_out[14]) );
    NR2 U100 ( .A(n298), .B(pop_empty), .Z(data_out[13]) );
    NR2 U101 ( .A(n299), .B(pop_empty), .Z(data_out[12]) );
    NR2 U102 ( .A(n300), .B(pop_empty), .Z(data_out[11]) );
    NR2 U103 ( .A(n301), .B(pop_empty), .Z(data_out[10]) );
    NR2 U104 ( .A(n302), .B(pop_empty), .Z(data_out[9]) );
    NR2 U105 ( .A(n303), .B(pop_empty), .Z(data_out[8]) );
    NR2 U106 ( .A(n304), .B(pop_empty), .Z(data_out[7]) );
    NR2 U107 ( .A(n305), .B(pop_empty), .Z(data_out[6]) );
    NR2 U108 ( .A(n306), .B(pop_empty), .Z(data_out[5]) );
    NR2 U109 ( .A(n307), .B(pop_empty), .Z(data_out[4]) );
    NR2 U110 ( .A(n308), .B(pop_empty), .Z(data_out[3]) );
    NR2 U111 ( .A(n309), .B(pop_empty), .Z(data_out[2]) );
    NR2 U112 ( .A(n310), .B(pop_empty), .Z(data_out[1]) );
    NR2 U113 ( .A(n311), .B(pop_empty), .Z(data_out[0]) );
    IV U114 ( .A(\dataout[9] ), .Z(n302) );
    IV U115 ( .A(\dataout[8] ), .Z(n303) );
    IV U116 ( .A(\dataout[7] ), .Z(n304) );
    IV U117 ( .A(\dataout[6] ), .Z(n305) );
    IV U118 ( .A(\dataout[5] ), .Z(n306) );
    IV U119 ( .A(\dataout[4] ), .Z(n307) );
    IV U120 ( .A(\dataout[3] ), .Z(n308) );
    IV U121 ( .A(\dataout[31] ), .Z(n280) );
    IV U122 ( .A(\dataout[30] ), .Z(n281) );
    IV U123 ( .A(\dataout[2] ), .Z(n309) );
    IV U124 ( .A(\dataout[29] ), .Z(n282) );
    IV U125 ( .A(\dataout[28] ), .Z(n283) );
    IV U126 ( .A(\dataout[27] ), .Z(n284) );
    IV U127 ( .A(\dataout[26] ), .Z(n285) );
    IV U128 ( .A(\dataout[25] ), .Z(n286) );
    IV U129 ( .A(\dataout[24] ), .Z(n287) );
    IV U130 ( .A(\dataout[23] ), .Z(n288) );
    IV U131 ( .A(\dataout[22] ), .Z(n289) );
    IV U132 ( .A(\dataout[21] ), .Z(n290) );
    IV U133 ( .A(\dataout[20] ), .Z(n291) );
    IV U134 ( .A(\dataout[1] ), .Z(n310) );
    IV U135 ( .A(\dataout[19] ), .Z(n292) );
    IV U136 ( .A(\dataout[18] ), .Z(n293) );
    IV U137 ( .A(\dataout[17] ), .Z(n294) );
    IV U138 ( .A(\dataout[16] ), .Z(n295) );
    IV U139 ( .A(\dataout[15] ), .Z(n296) );
    IV U140 ( .A(\dataout[14] ), .Z(n297) );
    IV U141 ( .A(\dataout[13] ), .Z(n298) );
    IV U142 ( .A(\dataout[12] ), .Z(n299) );
    IV U143 ( .A(\dataout[11] ), .Z(n300) );
    IV U144 ( .A(\dataout[10] ), .Z(n301) );
    IV U145 ( .A(\dataout[0] ), .Z(n311) );
endmodule

