// Write you SystemVerilog Assertions here !
